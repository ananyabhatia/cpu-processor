module wallacetree(A, B, O, overflow, ready, clk, ctrl_MULT);
   input [31:0] A, B;
   output [63:0] O;

    //full_adder(S, Cout, A, B, Cin);

    // A = y
    // B = x

    // wires with k are the output of the and gates
    wire k0_0, k0_1, k0_2, k0_3, k0_4, k0_5, k0_6, k0_7, k0_8, k0_9, k0_10, k0_11, k0_12, k0_13, k0_14, k0_15, k0_16, k0_17, k0_18, k0_19, k0_20, k0_21, k0_22, k0_23, k0_24, k0_25, k0_26, k0_27, k0_28, k0_29, k0_30, k0_31;

    assign k0_0  = A[0]  & B[0];
    assign k0_1  = A[0]  & B[1];
    assign k0_2  = A[0]  & B[2];
    assign k0_3  = A[0]  & B[3];
    assign k0_4  = A[0]  & B[4];
    assign k0_5  = A[0]  & B[5];
    assign k0_6  = A[0]  & B[6];
    assign k0_7  = A[0]  & B[7];
    assign k0_8  = A[0]  & B[8];
    assign k0_9  = A[0]  & B[9];
    assign k0_10 = A[0]  & B[10];
    assign k0_11 = A[0]  & B[11];
    assign k0_12 = A[0]  & B[12];
    assign k0_13 = A[0]  & B[13];
    assign k0_14 = A[0]  & B[14];
    assign k0_15 = A[0]  & B[15];
    assign k0_16 = A[0]  & B[16];
    assign k0_17 = A[0]  & B[17];
    assign k0_18 = A[0]  & B[18];
    assign k0_19 = A[0]  & B[19];
    assign k0_20 = A[0]  & B[20];
    assign k0_21 = A[0]  & B[21];
    assign k0_22 = A[0]  & B[22];
    assign k0_23 = A[0]  & B[23];
    assign k0_24 = A[0]  & B[24];
    assign k0_25 = A[0]  & B[25];
    assign k0_26 = A[0]  & B[26];
    assign k0_27 = A[0]  & B[27];
    assign k0_28 = A[0]  & B[28];
    assign k0_29 = A[0]  & B[29];
    assign k0_30 = A[0]  & B[30];
    assign k0_31 = !(A[0]  & B[31]);

    // Row 1
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k1_1;
    wire co11;
    full_adder adder11(k1_1, co11, k0_1, A[1] & B[0], 1'b0);
    wire k1_2;
    wire co12;
    full_adder adder12(k1_2, co12, k0_2, A[1] & B[1], co11);
    wire k1_3;
    wire co13;
    full_adder adder13(k1_3, co13, k0_3, A[1] & B[2], co12);
    wire k1_4;
    wire co14;
    full_adder adder14(k1_4, co14, k0_4, A[1] & B[3], co13);
    wire k1_5;
    wire co15;
    full_adder adder15(k1_5, co15, k0_5, A[1] & B[4], co14);
    wire k1_6;
    wire co16;
    full_adder adder16(k1_6, co16, k0_6, A[1] & B[5], co15);
    wire k1_7;
    wire co17;
    full_adder adder17(k1_7, co17, k0_7, A[1] & B[6], co16);
    wire k1_8;
    wire co18;
    full_adder adder18(k1_8, co18, k0_8, A[1] & B[7], co17);
    wire k1_9;
    wire co19;
    full_adder adder19(k1_9, co19, k0_9, A[1] & B[8], co18);
    wire k1_10;
    wire co110;
    full_adder adder110(k1_10, co110, k0_10, A[1] & B[9], co19);
    wire k1_11;
    wire co111;
    full_adder adder111(k1_11, co111, k0_11, A[1] & B[10], co110);
    wire k1_12;
    wire co112;
    full_adder adder112(k1_12, co112, k0_12, A[1] & B[11], co111);
    wire k1_13;
    wire co113;
    full_adder adder113(k1_13, co113, k0_13, A[1] & B[12], co112);
    wire k1_14;
    wire co114;
    full_adder adder114(k1_14, co114, k0_14, A[1] & B[13], co113);
    wire k1_15;
    wire co115;
    full_adder adder115(k1_15, co115, k0_15, A[1] & B[14], co114);
    wire k1_16;
    wire co116;
    full_adder adder116(k1_16, co116, k0_16, A[1] & B[15], co115);
    wire k1_17;
    wire co117;
    full_adder adder117(k1_17, co117, k0_17, A[1] & B[16], co116);
    wire k1_18;
    wire co118;
    full_adder adder118(k1_18, co118, k0_18, A[1] & B[17], co117);
    wire k1_19;
    wire co119;
    full_adder adder119(k1_19, co119, k0_19, A[1] & B[18], co118);
    wire k1_20;
    wire co120;
    full_adder adder120(k1_20, co120, k0_20, A[1] & B[19], co119);
    wire k1_21;
    wire co121;
    full_adder adder121(k1_21, co121, k0_21, A[1] & B[20], co120);
    wire k1_22;
    wire co122;
    full_adder adder122(k1_22, co122, k0_22, A[1] & B[21], co121);
    wire k1_23;
    wire co123;
    full_adder adder123(k1_23, co123, k0_23, A[1] & B[22], co122);
    wire k1_24;
    wire co124;
    full_adder adder124(k1_24, co124, k0_24, A[1] & B[23], co123);
    wire k1_25;
    wire co125;
    full_adder adder125(k1_25, co125, k0_25, A[1] & B[24], co124);
    wire k1_26;
    wire co126;
    full_adder adder126(k1_26, co126, k0_26, A[1] & B[25], co125);
    wire k1_27;
    wire co127;
    full_adder adder127(k1_27, co127, k0_27, A[1] & B[26], co126);
    wire k1_28;
    wire co128;
    full_adder adder128(k1_28, co128, k0_28, A[1] & B[27], co127);
    wire k1_29;
    wire co129;
    full_adder adder129(k1_29, co129, k0_29, A[1] & B[28], co128);
    wire k1_30;
    wire co130;
    full_adder adder130(k1_30, co130, k0_30, A[1] & B[29], co129);
    wire k1_31;
    wire co131;
    full_adder adder131(k1_31, co131, k0_31, A[1] & B[30], co130);
    wire k1_32;
    wire co132;
    full_adder adder132(k1_32, co132, 1'b1, !(A[1] & B[31]), co131);
    // Row 2
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k2_2;
    wire co22;
    full_adder adder22(k2_2, co22, k1_2, A[2] & B[0], 1'b0);
    wire k2_3;
    wire co23;
    full_adder adder23(k2_3, co23, k1_3, A[2] & B[1], co22);
    wire k2_4;
    wire co24;
    full_adder adder24(k2_4, co24, k1_4, A[2] & B[2], co23);
    wire k2_5;
    wire co25;
    full_adder adder25(k2_5, co25, k1_5, A[2] & B[3], co24);
    wire k2_6;
    wire co26;
    full_adder adder26(k2_6, co26, k1_6, A[2] & B[4], co25);
    wire k2_7;
    wire co27;
    full_adder adder27(k2_7, co27, k1_7, A[2] & B[5], co26);
    wire k2_8;
    wire co28;
    full_adder adder28(k2_8, co28, k1_8, A[2] & B[6], co27);
    wire k2_9;
    wire co29;
    full_adder adder29(k2_9, co29, k1_9, A[2] & B[7], co28);
    wire k2_10;
    wire co210;
    full_adder adder210(k2_10, co210, k1_10, A[2] & B[8], co29);
    wire k2_11;
    wire co211;
    full_adder adder211(k2_11, co211, k1_11, A[2] & B[9], co210);
    wire k2_12;
    wire co212;
    full_adder adder212(k2_12, co212, k1_12, A[2] & B[10], co211);
    wire k2_13;
    wire co213;
    full_adder adder213(k2_13, co213, k1_13, A[2] & B[11], co212);
    wire k2_14;
    wire co214;
    full_adder adder214(k2_14, co214, k1_14, A[2] & B[12], co213);
    wire k2_15;
    wire co215;
    full_adder adder215(k2_15, co215, k1_15, A[2] & B[13], co214);
    wire k2_16;
    wire co216;
    full_adder adder216(k2_16, co216, k1_16, A[2] & B[14], co215);
    wire k2_17;
    wire co217;
    full_adder adder217(k2_17, co217, k1_17, A[2] & B[15], co216);
    wire k2_18;
    wire co218;
    full_adder adder218(k2_18, co218, k1_18, A[2] & B[16], co217);
    wire k2_19;
    wire co219;
    full_adder adder219(k2_19, co219, k1_19, A[2] & B[17], co218);
    wire k2_20;
    wire co220;
    full_adder adder220(k2_20, co220, k1_20, A[2] & B[18], co219);
    wire k2_21;
    wire co221;
    full_adder adder221(k2_21, co221, k1_21, A[2] & B[19], co220);
    wire k2_22;
    wire co222;
    full_adder adder222(k2_22, co222, k1_22, A[2] & B[20], co221);
    wire k2_23;
    wire co223;
    full_adder adder223(k2_23, co223, k1_23, A[2] & B[21], co222);
    wire k2_24;
    wire co224;
    full_adder adder224(k2_24, co224, k1_24, A[2] & B[22], co223);
    wire k2_25;
    wire co225;
    full_adder adder225(k2_25, co225, k1_25, A[2] & B[23], co224);
    wire k2_26;
    wire co226;
    full_adder adder226(k2_26, co226, k1_26, A[2] & B[24], co225);
    wire k2_27;
    wire co227;
    full_adder adder227(k2_27, co227, k1_27, A[2] & B[25], co226);
    wire k2_28;
    wire co228;
    full_adder adder228(k2_28, co228, k1_28, A[2] & B[26], co227);
    wire k2_29;
    wire co229;
    full_adder adder229(k2_29, co229, k1_29, A[2] & B[27], co228);
    wire k2_30;
    wire co230;
    full_adder adder230(k2_30, co230, k1_30, A[2] & B[28], co229);
    wire k2_31;
    wire co231;
    full_adder adder231(k2_31, co231, k1_31, A[2] & B[29], co230);
    wire k2_32;
    wire co232;
    full_adder adder232(k2_32, co232, k1_32, A[2] & B[30], co231);
    wire k2_33;
    wire co233;
    full_adder adder233(k2_33, co233, co132, !(A[2] & B[31]), co232);
    // Row 3
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k3_3;
    wire co33;
    full_adder adder33(k3_3, co33, k2_3, A[3] & B[0], 1'b0);
    wire k3_4;
    wire co34;
    full_adder adder34(k3_4, co34, k2_4, A[3] & B[1], co33);
    wire k3_5;
    wire co35;
    full_adder adder35(k3_5, co35, k2_5, A[3] & B[2], co34);
    wire k3_6;
    wire co36;
    full_adder adder36(k3_6, co36, k2_6, A[3] & B[3], co35);
    wire k3_7;
    wire co37;
    full_adder adder37(k3_7, co37, k2_7, A[3] & B[4], co36);
    wire k3_8;
    wire co38;
    full_adder adder38(k3_8, co38, k2_8, A[3] & B[5], co37);
    wire k3_9;
    wire co39;
    full_adder adder39(k3_9, co39, k2_9, A[3] & B[6], co38);
    wire k3_10;
    wire co310;
    full_adder adder310(k3_10, co310, k2_10, A[3] & B[7], co39);
    wire k3_11;
    wire co311;
    full_adder adder311(k3_11, co311, k2_11, A[3] & B[8], co310);
    wire k3_12;
    wire co312;
    full_adder adder312(k3_12, co312, k2_12, A[3] & B[9], co311);
    wire k3_13;
    wire co313;
    full_adder adder313(k3_13, co313, k2_13, A[3] & B[10], co312);
    wire k3_14;
    wire co314;
    full_adder adder314(k3_14, co314, k2_14, A[3] & B[11], co313);
    wire k3_15;
    wire co315;
    full_adder adder315(k3_15, co315, k2_15, A[3] & B[12], co314);
    wire k3_16;
    wire co316;
    full_adder adder316(k3_16, co316, k2_16, A[3] & B[13], co315);
    wire k3_17;
    wire co317;
    full_adder adder317(k3_17, co317, k2_17, A[3] & B[14], co316);
    wire k3_18;
    wire co318;
    full_adder adder318(k3_18, co318, k2_18, A[3] & B[15], co317);
    wire k3_19;
    wire co319;
    full_adder adder319(k3_19, co319, k2_19, A[3] & B[16], co318);
    wire k3_20;
    wire co320;
    full_adder adder320(k3_20, co320, k2_20, A[3] & B[17], co319);
    wire k3_21;
    wire co321;
    full_adder adder321(k3_21, co321, k2_21, A[3] & B[18], co320);
    wire k3_22;
    wire co322;
    full_adder adder322(k3_22, co322, k2_22, A[3] & B[19], co321);
    wire k3_23;
    wire co323;
    full_adder adder323(k3_23, co323, k2_23, A[3] & B[20], co322);
    wire k3_24;
    wire co324;
    full_adder adder324(k3_24, co324, k2_24, A[3] & B[21], co323);
    wire k3_25;
    wire co325;
    full_adder adder325(k3_25, co325, k2_25, A[3] & B[22], co324);
    wire k3_26;
    wire co326;
    full_adder adder326(k3_26, co326, k2_26, A[3] & B[23], co325);
    wire k3_27;
    wire co327;
    full_adder adder327(k3_27, co327, k2_27, A[3] & B[24], co326);
    wire k3_28;
    wire co328;
    full_adder adder328(k3_28, co328, k2_28, A[3] & B[25], co327);
    wire k3_29;
    wire co329;
    full_adder adder329(k3_29, co329, k2_29, A[3] & B[26], co328);
    wire k3_30;
    wire co330;
    full_adder adder330(k3_30, co330, k2_30, A[3] & B[27], co329);
    wire k3_31;
    wire co331;
    full_adder adder331(k3_31, co331, k2_31, A[3] & B[28], co330);
    wire k3_32;
    wire co332;
    full_adder adder332(k3_32, co332, k2_32, A[3] & B[29], co331);
    wire k3_33;
    wire co333;
    full_adder adder333(k3_33, co333, k2_33, A[3] & B[30], co332);
    wire k3_34;
    wire co334;
    full_adder adder334(k3_34, co334, co233, !(A[3] & B[31]), co333);
    // Row 4
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k4_4;
    wire co44;
    full_adder adder44(k4_4, co44, k3_4, A[4] & B[0], 1'b0);
    wire k4_5;
    wire co45;
    full_adder adder45(k4_5, co45, k3_5, A[4] & B[1], co44);
    wire k4_6;
    wire co46;
    full_adder adder46(k4_6, co46, k3_6, A[4] & B[2], co45);
    wire k4_7;
    wire co47;
    full_adder adder47(k4_7, co47, k3_7, A[4] & B[3], co46);
    wire k4_8;
    wire co48;
    full_adder adder48(k4_8, co48, k3_8, A[4] & B[4], co47);
    wire k4_9;
    wire co49;
    full_adder adder49(k4_9, co49, k3_9, A[4] & B[5], co48);
    wire k4_10;
    wire co410;
    full_adder adder410(k4_10, co410, k3_10, A[4] & B[6], co49);
    wire k4_11;
    wire co411;
    full_adder adder411(k4_11, co411, k3_11, A[4] & B[7], co410);
    wire k4_12;
    wire co412;
    full_adder adder412(k4_12, co412, k3_12, A[4] & B[8], co411);
    wire k4_13;
    wire co413;
    full_adder adder413(k4_13, co413, k3_13, A[4] & B[9], co412);
    wire k4_14;
    wire co414;
    full_adder adder414(k4_14, co414, k3_14, A[4] & B[10], co413);
    wire k4_15;
    wire co415;
    full_adder adder415(k4_15, co415, k3_15, A[4] & B[11], co414);
    wire k4_16;
    wire co416;
    full_adder adder416(k4_16, co416, k3_16, A[4] & B[12], co415);
    wire k4_17;
    wire co417;
    full_adder adder417(k4_17, co417, k3_17, A[4] & B[13], co416);
    wire k4_18;
    wire co418;
    full_adder adder418(k4_18, co418, k3_18, A[4] & B[14], co417);
    wire k4_19;
    wire co419;
    full_adder adder419(k4_19, co419, k3_19, A[4] & B[15], co418);
    wire k4_20;
    wire co420;
    full_adder adder420(k4_20, co420, k3_20, A[4] & B[16], co419);
    wire k4_21;
    wire co421;
    full_adder adder421(k4_21, co421, k3_21, A[4] & B[17], co420);
    wire k4_22;
    wire co422;
    full_adder adder422(k4_22, co422, k3_22, A[4] & B[18], co421);
    wire k4_23;
    wire co423;
    full_adder adder423(k4_23, co423, k3_23, A[4] & B[19], co422);
    wire k4_24;
    wire co424;
    full_adder adder424(k4_24, co424, k3_24, A[4] & B[20], co423);
    wire k4_25;
    wire co425;
    full_adder adder425(k4_25, co425, k3_25, A[4] & B[21], co424);
    wire k4_26;
    wire co426;
    full_adder adder426(k4_26, co426, k3_26, A[4] & B[22], co425);
    wire k4_27;
    wire co427;
    full_adder adder427(k4_27, co427, k3_27, A[4] & B[23], co426);
    wire k4_28;
    wire co428;
    full_adder adder428(k4_28, co428, k3_28, A[4] & B[24], co427);
    wire k4_29;
    wire co429;
    full_adder adder429(k4_29, co429, k3_29, A[4] & B[25], co428);
    wire k4_30;
    wire co430;
    full_adder adder430(k4_30, co430, k3_30, A[4] & B[26], co429);
    wire k4_31;
    wire co431;
    full_adder adder431(k4_31, co431, k3_31, A[4] & B[27], co430);
    wire k4_32;
    wire co432;
    full_adder adder432(k4_32, co432, k3_32, A[4] & B[28], co431);
    wire k4_33;
    wire co433;
    full_adder adder433(k4_33, co433, k3_33, A[4] & B[29], co432);
    wire k4_34;
    wire co434;
    full_adder adder434(k4_34, co434, k3_34, A[4] & B[30], co433);
    wire k4_35;
    wire co435;
    full_adder adder435(k4_35, co435, co334, !(A[4] & B[31]), co434);
    // Row 5
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k5_5;
    wire co55;
    full_adder adder55(k5_5, co55, k4_5, A[5] & B[0], 1'b0);
    wire k5_6;
    wire co56;
    full_adder adder56(k5_6, co56, k4_6, A[5] & B[1], co55);
    wire k5_7;
    wire co57;
    full_adder adder57(k5_7, co57, k4_7, A[5] & B[2], co56);
    wire k5_8;
    wire co58;
    full_adder adder58(k5_8, co58, k4_8, A[5] & B[3], co57);
    wire k5_9;
    wire co59;
    full_adder adder59(k5_9, co59, k4_9, A[5] & B[4], co58);
    wire k5_10;
    wire co510;
    full_adder adder510(k5_10, co510, k4_10, A[5] & B[5], co59);
    wire k5_11;
    wire co511;
    full_adder adder511(k5_11, co511, k4_11, A[5] & B[6], co510);
    wire k5_12;
    wire co512;
    full_adder adder512(k5_12, co512, k4_12, A[5] & B[7], co511);
    wire k5_13;
    wire co513;
    full_adder adder513(k5_13, co513, k4_13, A[5] & B[8], co512);
    wire k5_14;
    wire co514;
    full_adder adder514(k5_14, co514, k4_14, A[5] & B[9], co513);
    wire k5_15;
    wire co515;
    full_adder adder515(k5_15, co515, k4_15, A[5] & B[10], co514);
    wire k5_16;
    wire co516;
    full_adder adder516(k5_16, co516, k4_16, A[5] & B[11], co515);
    wire k5_17;
    wire co517;
    full_adder adder517(k5_17, co517, k4_17, A[5] & B[12], co516);
    wire k5_18;
    wire co518;
    full_adder adder518(k5_18, co518, k4_18, A[5] & B[13], co517);
    wire k5_19;
    wire co519;
    full_adder adder519(k5_19, co519, k4_19, A[5] & B[14], co518);
    wire k5_20;
    wire co520;
    full_adder adder520(k5_20, co520, k4_20, A[5] & B[15], co519);
    wire k5_21;
    wire co521;
    full_adder adder521(k5_21, co521, k4_21, A[5] & B[16], co520);
    wire k5_22;
    wire co522;
    full_adder adder522(k5_22, co522, k4_22, A[5] & B[17], co521);
    wire k5_23;
    wire co523;
    full_adder adder523(k5_23, co523, k4_23, A[5] & B[18], co522);
    wire k5_24;
    wire co524;
    full_adder adder524(k5_24, co524, k4_24, A[5] & B[19], co523);
    wire k5_25;
    wire co525;
    full_adder adder525(k5_25, co525, k4_25, A[5] & B[20], co524);
    wire k5_26;
    wire co526;
    full_adder adder526(k5_26, co526, k4_26, A[5] & B[21], co525);
    wire k5_27;
    wire co527;
    full_adder adder527(k5_27, co527, k4_27, A[5] & B[22], co526);
    wire k5_28;
    wire co528;
    full_adder adder528(k5_28, co528, k4_28, A[5] & B[23], co527);
    wire k5_29;
    wire co529;
    full_adder adder529(k5_29, co529, k4_29, A[5] & B[24], co528);
    wire k5_30;
    wire co530;
    full_adder adder530(k5_30, co530, k4_30, A[5] & B[25], co529);
    wire k5_31;
    wire co531;
    full_adder adder531(k5_31, co531, k4_31, A[5] & B[26], co530);
    wire k5_32;
    wire co532;
    full_adder adder532(k5_32, co532, k4_32, A[5] & B[27], co531);
    wire k5_33;
    wire co533;
    full_adder adder533(k5_33, co533, k4_33, A[5] & B[28], co532);
    wire k5_34;
    wire co534;
    full_adder adder534(k5_34, co534, k4_34, A[5] & B[29], co533);
    wire k5_35;
    wire co535;
    full_adder adder535(k5_35, co535, k4_35, A[5] & B[30], co534);
    wire k5_36;
    wire co536;
    full_adder adder536(k5_36, co536, co435, !(A[5] & B[31]), co535);
    // Row 6
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k6_6;
    wire co66;
    full_adder adder66(k6_6, co66, k5_6, A[6] & B[0], 1'b0);
    wire k6_7;
    wire co67;
    full_adder adder67(k6_7, co67, k5_7, A[6] & B[1], co66);
    wire k6_8;
    wire co68;
    full_adder adder68(k6_8, co68, k5_8, A[6] & B[2], co67);
    wire k6_9;
    wire co69;
    full_adder adder69(k6_9, co69, k5_9, A[6] & B[3], co68);
    wire k6_10;
    wire co610;
    full_adder adder610(k6_10, co610, k5_10, A[6] & B[4], co69);
    wire k6_11;
    wire co611;
    full_adder adder611(k6_11, co611, k5_11, A[6] & B[5], co610);
    wire k6_12;
    wire co612;
    full_adder adder612(k6_12, co612, k5_12, A[6] & B[6], co611);
    wire k6_13;
    wire co613;
    full_adder adder613(k6_13, co613, k5_13, A[6] & B[7], co612);
    wire k6_14;
    wire co614;
    full_adder adder614(k6_14, co614, k5_14, A[6] & B[8], co613);
    wire k6_15;
    wire co615;
    full_adder adder615(k6_15, co615, k5_15, A[6] & B[9], co614);
    wire k6_16;
    wire co616;
    full_adder adder616(k6_16, co616, k5_16, A[6] & B[10], co615);
    wire k6_17;
    wire co617;
    full_adder adder617(k6_17, co617, k5_17, A[6] & B[11], co616);
    wire k6_18;
    wire co618;
    full_adder adder618(k6_18, co618, k5_18, A[6] & B[12], co617);
    wire k6_19;
    wire co619;
    full_adder adder619(k6_19, co619, k5_19, A[6] & B[13], co618);
    wire k6_20;
    wire co620;
    full_adder adder620(k6_20, co620, k5_20, A[6] & B[14], co619);
    wire k6_21;
    wire co621;
    full_adder adder621(k6_21, co621, k5_21, A[6] & B[15], co620);
    wire k6_22;
    wire co622;
    full_adder adder622(k6_22, co622, k5_22, A[6] & B[16], co621);
    wire k6_23;
    wire co623;
    full_adder adder623(k6_23, co623, k5_23, A[6] & B[17], co622);
    wire k6_24;
    wire co624;
    full_adder adder624(k6_24, co624, k5_24, A[6] & B[18], co623);
    wire k6_25;
    wire co625;
    full_adder adder625(k6_25, co625, k5_25, A[6] & B[19], co624);
    wire k6_26;
    wire co626;
    full_adder adder626(k6_26, co626, k5_26, A[6] & B[20], co625);
    wire k6_27;
    wire co627;
    full_adder adder627(k6_27, co627, k5_27, A[6] & B[21], co626);
    wire k6_28;
    wire co628;
    full_adder adder628(k6_28, co628, k5_28, A[6] & B[22], co627);
    wire k6_29;
    wire co629;
    full_adder adder629(k6_29, co629, k5_29, A[6] & B[23], co628);
    wire k6_30;
    wire co630;
    full_adder adder630(k6_30, co630, k5_30, A[6] & B[24], co629);
    wire k6_31;
    wire co631;
    full_adder adder631(k6_31, co631, k5_31, A[6] & B[25], co630);
    wire k6_32;
    wire co632;
    full_adder adder632(k6_32, co632, k5_32, A[6] & B[26], co631);
    wire k6_33;
    wire co633;
    full_adder adder633(k6_33, co633, k5_33, A[6] & B[27], co632);
    wire k6_34;
    wire co634;
    full_adder adder634(k6_34, co634, k5_34, A[6] & B[28], co633);
    wire k6_35;
    wire co635;
    full_adder adder635(k6_35, co635, k5_35, A[6] & B[29], co634);
    wire k6_36;
    wire co636;
    full_adder adder636(k6_36, co636, k5_36, A[6] & B[30], co635);
    wire k6_37;
    wire co637;
    full_adder adder637(k6_37, co637, co536, !(A[6] & B[31]), co636);
    // Row 7
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k7_7;
    wire co77;
    full_adder adder77(k7_7, co77, k6_7, A[7] & B[0], 1'b0);
    wire k7_8;
    wire co78;
    full_adder adder78(k7_8, co78, k6_8, A[7] & B[1], co77);
    wire k7_9;
    wire co79;
    full_adder adder79(k7_9, co79, k6_9, A[7] & B[2], co78);
    wire k7_10;
    wire co710;
    full_adder adder710(k7_10, co710, k6_10, A[7] & B[3], co79);
    wire k7_11;
    wire co711;
    full_adder adder711(k7_11, co711, k6_11, A[7] & B[4], co710);
    wire k7_12;
    wire co712;
    full_adder adder712(k7_12, co712, k6_12, A[7] & B[5], co711);
    wire k7_13;
    wire co713;
    full_adder adder713(k7_13, co713, k6_13, A[7] & B[6], co712);
    wire k7_14;
    wire co714;
    full_adder adder714(k7_14, co714, k6_14, A[7] & B[7], co713);
    wire k7_15;
    wire co715;
    full_adder adder715(k7_15, co715, k6_15, A[7] & B[8], co714);
    wire k7_16;
    wire co716;
    full_adder adder716(k7_16, co716, k6_16, A[7] & B[9], co715);
    wire k7_17;
    wire co717;
    full_adder adder717(k7_17, co717, k6_17, A[7] & B[10], co716);
    wire k7_18;
    wire co718;
    full_adder adder718(k7_18, co718, k6_18, A[7] & B[11], co717);
    wire k7_19;
    wire co719;
    full_adder adder719(k7_19, co719, k6_19, A[7] & B[12], co718);
    wire k7_20;
    wire co720;
    full_adder adder720(k7_20, co720, k6_20, A[7] & B[13], co719);
    wire k7_21;
    wire co721;
    full_adder adder721(k7_21, co721, k6_21, A[7] & B[14], co720);
    wire k7_22;
    wire co722;
    full_adder adder722(k7_22, co722, k6_22, A[7] & B[15], co721);
    wire k7_23;
    wire co723;
    full_adder adder723(k7_23, co723, k6_23, A[7] & B[16], co722);
    wire k7_24;
    wire co724;
    full_adder adder724(k7_24, co724, k6_24, A[7] & B[17], co723);
    wire k7_25;
    wire co725;
    full_adder adder725(k7_25, co725, k6_25, A[7] & B[18], co724);
    wire k7_26;
    wire co726;
    full_adder adder726(k7_26, co726, k6_26, A[7] & B[19], co725);
    wire k7_27;
    wire co727;
    full_adder adder727(k7_27, co727, k6_27, A[7] & B[20], co726);
    wire k7_28;
    wire co728;
    full_adder adder728(k7_28, co728, k6_28, A[7] & B[21], co727);
    wire k7_29;
    wire co729;
    full_adder adder729(k7_29, co729, k6_29, A[7] & B[22], co728);
    wire k7_30;
    wire co730;
    full_adder adder730(k7_30, co730, k6_30, A[7] & B[23], co729);
    wire k7_31;
    wire co731;
    full_adder adder731(k7_31, co731, k6_31, A[7] & B[24], co730);
    wire k7_32;
    wire co732;
    full_adder adder732(k7_32, co732, k6_32, A[7] & B[25], co731);
    wire k7_33;
    wire co733;
    full_adder adder733(k7_33, co733, k6_33, A[7] & B[26], co732);
    wire k7_34;
    wire co734;
    full_adder adder734(k7_34, co734, k6_34, A[7] & B[27], co733);
    wire k7_35;
    wire co735;
    full_adder adder735(k7_35, co735, k6_35, A[7] & B[28], co734);
    wire k7_36;
    wire co736;
    full_adder adder736(k7_36, co736, k6_36, A[7] & B[29], co735);
    wire k7_37;
    wire co737;
    full_adder adder737(k7_37, co737, k6_37, A[7] & B[30], co736);
    wire k7_38;
    wire co738;
    full_adder adder738(k7_38, co738, co637, !(A[7] & B[31]), co737);
    // Row 8
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k8_8;
    wire co88;
    full_adder adder88(k8_8, co88, k7_8, A[8] & B[0], 1'b0);
    wire k8_9;
    wire co89;
    full_adder adder89(k8_9, co89, k7_9, A[8] & B[1], co88);
    wire k8_10;
    wire co810;
    full_adder adder810(k8_10, co810, k7_10, A[8] & B[2], co89);
    wire k8_11;
    wire co811;
    full_adder adder811(k8_11, co811, k7_11, A[8] & B[3], co810);
    wire k8_12;
    wire co812;
    full_adder adder812(k8_12, co812, k7_12, A[8] & B[4], co811);
    wire k8_13;
    wire co813;
    full_adder adder813(k8_13, co813, k7_13, A[8] & B[5], co812);
    wire k8_14;
    wire co814;
    full_adder adder814(k8_14, co814, k7_14, A[8] & B[6], co813);
    wire k8_15;
    wire co815;
    full_adder adder815(k8_15, co815, k7_15, A[8] & B[7], co814);
    wire k8_16;
    wire co816;
    full_adder adder816(k8_16, co816, k7_16, A[8] & B[8], co815);
    wire k8_17;
    wire co817;
    full_adder adder817(k8_17, co817, k7_17, A[8] & B[9], co816);
    wire k8_18;
    wire co818;
    full_adder adder818(k8_18, co818, k7_18, A[8] & B[10], co817);
    wire k8_19;
    wire co819;
    full_adder adder819(k8_19, co819, k7_19, A[8] & B[11], co818);
    wire k8_20;
    wire co820;
    full_adder adder820(k8_20, co820, k7_20, A[8] & B[12], co819);
    wire k8_21;
    wire co821;
    full_adder adder821(k8_21, co821, k7_21, A[8] & B[13], co820);
    wire k8_22;
    wire co822;
    full_adder adder822(k8_22, co822, k7_22, A[8] & B[14], co821);
    wire k8_23;
    wire co823;
    full_adder adder823(k8_23, co823, k7_23, A[8] & B[15], co822);
    wire k8_24;
    wire co824;
    full_adder adder824(k8_24, co824, k7_24, A[8] & B[16], co823);
    wire k8_25;
    wire co825;
    full_adder adder825(k8_25, co825, k7_25, A[8] & B[17], co824);
    wire k8_26;
    wire co826;
    full_adder adder826(k8_26, co826, k7_26, A[8] & B[18], co825);
    wire k8_27;
    wire co827;
    full_adder adder827(k8_27, co827, k7_27, A[8] & B[19], co826);
    wire k8_28;
    wire co828;
    full_adder adder828(k8_28, co828, k7_28, A[8] & B[20], co827);
    wire k8_29;
    wire co829;
    full_adder adder829(k8_29, co829, k7_29, A[8] & B[21], co828);
    wire k8_30;
    wire co830;
    full_adder adder830(k8_30, co830, k7_30, A[8] & B[22], co829);
    wire k8_31;
    wire co831;
    full_adder adder831(k8_31, co831, k7_31, A[8] & B[23], co830);
    wire k8_32;
    wire co832;
    full_adder adder832(k8_32, co832, k7_32, A[8] & B[24], co831);
    wire k8_33;
    wire co833;
    full_adder adder833(k8_33, co833, k7_33, A[8] & B[25], co832);
    wire k8_34;
    wire co834;
    full_adder adder834(k8_34, co834, k7_34, A[8] & B[26], co833);
    wire k8_35;
    wire co835;
    full_adder adder835(k8_35, co835, k7_35, A[8] & B[27], co834);
    wire k8_36;
    wire co836;
    full_adder adder836(k8_36, co836, k7_36, A[8] & B[28], co835);
    wire k8_37;
    wire co837;
    full_adder adder837(k8_37, co837, k7_37, A[8] & B[29], co836);
    wire k8_38;
    wire co838;
    full_adder adder838(k8_38, co838, k7_38, A[8] & B[30], co837);
    wire k8_39;
    wire co839;
    full_adder adder839(k8_39, co839, co738, !(A[8] & B[31]), co838);
    // Row 9
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k9_9;
    wire co99;
    full_adder adder99(k9_9, co99, k8_9, A[9] & B[0], 1'b0);
    wire k9_10;
    wire co910;
    full_adder adder910(k9_10, co910, k8_10, A[9] & B[1], co99);
    wire k9_11;
    wire co911;
    full_adder adder911(k9_11, co911, k8_11, A[9] & B[2], co910);
    wire k9_12;
    wire co912;
    full_adder adder912(k9_12, co912, k8_12, A[9] & B[3], co911);
    wire k9_13;
    wire co913;
    full_adder adder913(k9_13, co913, k8_13, A[9] & B[4], co912);
    wire k9_14;
    wire co914;
    full_adder adder914(k9_14, co914, k8_14, A[9] & B[5], co913);
    wire k9_15;
    wire co915;
    full_adder adder915(k9_15, co915, k8_15, A[9] & B[6], co914);
    wire k9_16;
    wire co916;
    full_adder adder916(k9_16, co916, k8_16, A[9] & B[7], co915);
    wire k9_17;
    wire co917;
    full_adder adder917(k9_17, co917, k8_17, A[9] & B[8], co916);
    wire k9_18;
    wire co918;
    full_adder adder918(k9_18, co918, k8_18, A[9] & B[9], co917);
    wire k9_19;
    wire co919;
    full_adder adder919(k9_19, co919, k8_19, A[9] & B[10], co918);
    wire k9_20;
    wire co920;
    full_adder adder920(k9_20, co920, k8_20, A[9] & B[11], co919);
    wire k9_21;
    wire co921;
    full_adder adder921(k9_21, co921, k8_21, A[9] & B[12], co920);
    wire k9_22;
    wire co922;
    full_adder adder922(k9_22, co922, k8_22, A[9] & B[13], co921);
    wire k9_23;
    wire co923;
    full_adder adder923(k9_23, co923, k8_23, A[9] & B[14], co922);
    wire k9_24;
    wire co924;
    full_adder adder924(k9_24, co924, k8_24, A[9] & B[15], co923);
    wire k9_25;
    wire co925;
    full_adder adder925(k9_25, co925, k8_25, A[9] & B[16], co924);
    wire k9_26;
    wire co926;
    full_adder adder926(k9_26, co926, k8_26, A[9] & B[17], co925);
    wire k9_27;
    wire co927;
    full_adder adder927(k9_27, co927, k8_27, A[9] & B[18], co926);
    wire k9_28;
    wire co928;
    full_adder adder928(k9_28, co928, k8_28, A[9] & B[19], co927);
    wire k9_29;
    wire co929;
    full_adder adder929(k9_29, co929, k8_29, A[9] & B[20], co928);
    wire k9_30;
    wire co930;
    full_adder adder930(k9_30, co930, k8_30, A[9] & B[21], co929);
    wire k9_31;
    wire co931;
    full_adder adder931(k9_31, co931, k8_31, A[9] & B[22], co930);
    wire k9_32;
    wire co932;
    full_adder adder932(k9_32, co932, k8_32, A[9] & B[23], co931);
    wire k9_33;
    wire co933;
    full_adder adder933(k9_33, co933, k8_33, A[9] & B[24], co932);
    wire k9_34;
    wire co934;
    full_adder adder934(k9_34, co934, k8_34, A[9] & B[25], co933);
    wire k9_35;
    wire co935;
    full_adder adder935(k9_35, co935, k8_35, A[9] & B[26], co934);
    wire k9_36;
    wire co936;
    full_adder adder936(k9_36, co936, k8_36, A[9] & B[27], co935);
    wire k9_37;
    wire co937;
    full_adder adder937(k9_37, co937, k8_37, A[9] & B[28], co936);
    wire k9_38;
    wire co938;
    full_adder adder938(k9_38, co938, k8_38, A[9] & B[29], co937);
    wire k9_39;
    wire co939;
    full_adder adder939(k9_39, co939, k8_39, A[9] & B[30], co938);
    wire k9_40;
    wire co940;
    full_adder adder940(k9_40, co940, co839, !(A[9] & B[31]), co939);
    // Row 10
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k10_10;
    wire co1010;
    full_adder adder1010(k10_10, co1010, k9_10, A[10] & B[0], 1'b0);
    wire k10_11;
    wire co1011;
    full_adder adder1011(k10_11, co1011, k9_11, A[10] & B[1], co1010);
    wire k10_12;
    wire co1012;
    full_adder adder1012(k10_12, co1012, k9_12, A[10] & B[2], co1011);
    wire k10_13;
    wire co1013;
    full_adder adder1013(k10_13, co1013, k9_13, A[10] & B[3], co1012);
    wire k10_14;
    wire co1014;
    full_adder adder1014(k10_14, co1014, k9_14, A[10] & B[4], co1013);
    wire k10_15;
    wire co1015;
    full_adder adder1015(k10_15, co1015, k9_15, A[10] & B[5], co1014);
    wire k10_16;
    wire co1016;
    full_adder adder1016(k10_16, co1016, k9_16, A[10] & B[6], co1015);
    wire k10_17;
    wire co1017;
    full_adder adder1017(k10_17, co1017, k9_17, A[10] & B[7], co1016);
    wire k10_18;
    wire co1018;
    full_adder adder1018(k10_18, co1018, k9_18, A[10] & B[8], co1017);
    wire k10_19;
    wire co1019;
    full_adder adder1019(k10_19, co1019, k9_19, A[10] & B[9], co1018);
    wire k10_20;
    wire co1020;
    full_adder adder1020(k10_20, co1020, k9_20, A[10] & B[10], co1019);
    wire k10_21;
    wire co1021;
    full_adder adder1021(k10_21, co1021, k9_21, A[10] & B[11], co1020);
    wire k10_22;
    wire co1022;
    full_adder adder1022(k10_22, co1022, k9_22, A[10] & B[12], co1021);
    wire k10_23;
    wire co1023;
    full_adder adder1023(k10_23, co1023, k9_23, A[10] & B[13], co1022);
    wire k10_24;
    wire co1024;
    full_adder adder1024(k10_24, co1024, k9_24, A[10] & B[14], co1023);
    wire k10_25;
    wire co1025;
    full_adder adder1025(k10_25, co1025, k9_25, A[10] & B[15], co1024);
    wire k10_26;
    wire co1026;
    full_adder adder1026(k10_26, co1026, k9_26, A[10] & B[16], co1025);
    wire k10_27;
    wire co1027;
    full_adder adder1027(k10_27, co1027, k9_27, A[10] & B[17], co1026);
    wire k10_28;
    wire co1028;
    full_adder adder1028(k10_28, co1028, k9_28, A[10] & B[18], co1027);
    wire k10_29;
    wire co1029;
    full_adder adder1029(k10_29, co1029, k9_29, A[10] & B[19], co1028);
    wire k10_30;
    wire co1030;
    full_adder adder1030(k10_30, co1030, k9_30, A[10] & B[20], co1029);
    wire k10_31;
    wire co1031;
    full_adder adder1031(k10_31, co1031, k9_31, A[10] & B[21], co1030);
    wire k10_32;
    wire co1032;
    full_adder adder1032(k10_32, co1032, k9_32, A[10] & B[22], co1031);
    wire k10_33;
    wire co1033;
    full_adder adder1033(k10_33, co1033, k9_33, A[10] & B[23], co1032);
    wire k10_34;
    wire co1034;
    full_adder adder1034(k10_34, co1034, k9_34, A[10] & B[24], co1033);
    wire k10_35;
    wire co1035;
    full_adder adder1035(k10_35, co1035, k9_35, A[10] & B[25], co1034);
    wire k10_36;
    wire co1036;
    full_adder adder1036(k10_36, co1036, k9_36, A[10] & B[26], co1035);
    wire k10_37;
    wire co1037;
    full_adder adder1037(k10_37, co1037, k9_37, A[10] & B[27], co1036);
    wire k10_38;
    wire co1038;
    full_adder adder1038(k10_38, co1038, k9_38, A[10] & B[28], co1037);
    wire k10_39;
    wire co1039;
    full_adder adder1039(k10_39, co1039, k9_39, A[10] & B[29], co1038);
    wire k10_40;
    wire co1040;
    full_adder adder1040(k10_40, co1040, k9_40, A[10] & B[30], co1039);
    wire k10_41;
    wire co1041;
    full_adder adder1041(k10_41, co1041, co940, !(A[10] & B[31]), co1040);
    // Row 11
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k11_11;
    wire co1111;
    full_adder adder1111(k11_11, co1111, k10_11, A[11] & B[0], 1'b0);
    wire k11_12;
    wire co1112;
    full_adder adder1112(k11_12, co1112, k10_12, A[11] & B[1], co1111);
    wire k11_13;
    wire co1113;
    full_adder adder1113(k11_13, co1113, k10_13, A[11] & B[2], co1112);
    wire k11_14;
    wire co1114;
    full_adder adder1114(k11_14, co1114, k10_14, A[11] & B[3], co1113);
    wire k11_15;
    wire co1115;
    full_adder adder1115(k11_15, co1115, k10_15, A[11] & B[4], co1114);
    wire k11_16;
    wire co1116;
    full_adder adder1116(k11_16, co1116, k10_16, A[11] & B[5], co1115);
    wire k11_17;
    wire co1117;
    full_adder adder1117(k11_17, co1117, k10_17, A[11] & B[6], co1116);
    wire k11_18;
    wire co1118;
    full_adder adder1118(k11_18, co1118, k10_18, A[11] & B[7], co1117);
    wire k11_19;
    wire co1119;
    full_adder adder1119(k11_19, co1119, k10_19, A[11] & B[8], co1118);
    wire k11_20;
    wire co1120;
    full_adder adder1120(k11_20, co1120, k10_20, A[11] & B[9], co1119);
    wire k11_21;
    wire co1121;
    full_adder adder1121(k11_21, co1121, k10_21, A[11] & B[10], co1120);
    wire k11_22;
    wire co1122;
    full_adder adder1122(k11_22, co1122, k10_22, A[11] & B[11], co1121);
    wire k11_23;
    wire co1123;
    full_adder adder1123(k11_23, co1123, k10_23, A[11] & B[12], co1122);
    wire k11_24;
    wire co1124;
    full_adder adder1124(k11_24, co1124, k10_24, A[11] & B[13], co1123);
    wire k11_25;
    wire co1125;
    full_adder adder1125(k11_25, co1125, k10_25, A[11] & B[14], co1124);
    wire k11_26;
    wire co1126;
    full_adder adder1126(k11_26, co1126, k10_26, A[11] & B[15], co1125);
    wire k11_27;
    wire co1127;
    full_adder adder1127(k11_27, co1127, k10_27, A[11] & B[16], co1126);
    wire k11_28;
    wire co1128;
    full_adder adder1128(k11_28, co1128, k10_28, A[11] & B[17], co1127);
    wire k11_29;
    wire co1129;
    full_adder adder1129(k11_29, co1129, k10_29, A[11] & B[18], co1128);
    wire k11_30;
    wire co1130;
    full_adder adder1130(k11_30, co1130, k10_30, A[11] & B[19], co1129);
    wire k11_31;
    wire co1131;
    full_adder adder1131(k11_31, co1131, k10_31, A[11] & B[20], co1130);
    wire k11_32;
    wire co1132;
    full_adder adder1132(k11_32, co1132, k10_32, A[11] & B[21], co1131);
    wire k11_33;
    wire co1133;
    full_adder adder1133(k11_33, co1133, k10_33, A[11] & B[22], co1132);
    wire k11_34;
    wire co1134;
    full_adder adder1134(k11_34, co1134, k10_34, A[11] & B[23], co1133);
    wire k11_35;
    wire co1135;
    full_adder adder1135(k11_35, co1135, k10_35, A[11] & B[24], co1134);
    wire k11_36;
    wire co1136;
    full_adder adder1136(k11_36, co1136, k10_36, A[11] & B[25], co1135);
    wire k11_37;
    wire co1137;
    full_adder adder1137(k11_37, co1137, k10_37, A[11] & B[26], co1136);
    wire k11_38;
    wire co1138;
    full_adder adder1138(k11_38, co1138, k10_38, A[11] & B[27], co1137);
    wire k11_39;
    wire co1139;
    full_adder adder1139(k11_39, co1139, k10_39, A[11] & B[28], co1138);
    wire k11_40;
    wire co1140;
    full_adder adder1140(k11_40, co1140, k10_40, A[11] & B[29], co1139);
    wire k11_41;
    wire co1141;
    full_adder adder1141(k11_41, co1141, k10_41, A[11] & B[30], co1140);
    wire k11_42;
    wire co1142;
    full_adder adder1142(k11_42, co1142, co1041, !(A[11] & B[31]), co1141);
    // Row 12
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k12_12;
    wire co1212;
    full_adder adder1212(k12_12, co1212, k11_12, A[12] & B[0], 1'b0);
    wire k12_13;
    wire co1213;
    full_adder adder1213(k12_13, co1213, k11_13, A[12] & B[1], co1212);
    wire k12_14;
    wire co1214;
    full_adder adder1214(k12_14, co1214, k11_14, A[12] & B[2], co1213);
    wire k12_15;
    wire co1215;
    full_adder adder1215(k12_15, co1215, k11_15, A[12] & B[3], co1214);
    wire k12_16;
    wire co1216;
    full_adder adder1216(k12_16, co1216, k11_16, A[12] & B[4], co1215);
    wire k12_17;
    wire co1217;
    full_adder adder1217(k12_17, co1217, k11_17, A[12] & B[5], co1216);
    wire k12_18;
    wire co1218;
    full_adder adder1218(k12_18, co1218, k11_18, A[12] & B[6], co1217);
    wire k12_19;
    wire co1219;
    full_adder adder1219(k12_19, co1219, k11_19, A[12] & B[7], co1218);
    wire k12_20;
    wire co1220;
    full_adder adder1220(k12_20, co1220, k11_20, A[12] & B[8], co1219);
    wire k12_21;
    wire co1221;
    full_adder adder1221(k12_21, co1221, k11_21, A[12] & B[9], co1220);
    wire k12_22;
    wire co1222;
    full_adder adder1222(k12_22, co1222, k11_22, A[12] & B[10], co1221);
    wire k12_23;
    wire co1223;
    full_adder adder1223(k12_23, co1223, k11_23, A[12] & B[11], co1222);
    wire k12_24;
    wire co1224;
    full_adder adder1224(k12_24, co1224, k11_24, A[12] & B[12], co1223);
    wire k12_25;
    wire co1225;
    full_adder adder1225(k12_25, co1225, k11_25, A[12] & B[13], co1224);
    wire k12_26;
    wire co1226;
    full_adder adder1226(k12_26, co1226, k11_26, A[12] & B[14], co1225);
    wire k12_27;
    wire co1227;
    full_adder adder1227(k12_27, co1227, k11_27, A[12] & B[15], co1226);
    wire k12_28;
    wire co1228;
    full_adder adder1228(k12_28, co1228, k11_28, A[12] & B[16], co1227);
    wire k12_29;
    wire co1229;
    full_adder adder1229(k12_29, co1229, k11_29, A[12] & B[17], co1228);
    wire k12_30;
    wire co1230;
    full_adder adder1230(k12_30, co1230, k11_30, A[12] & B[18], co1229);
    wire k12_31;
    wire co1231;
    full_adder adder1231(k12_31, co1231, k11_31, A[12] & B[19], co1230);
    wire k12_32;
    wire co1232;
    full_adder adder1232(k12_32, co1232, k11_32, A[12] & B[20], co1231);
    wire k12_33;
    wire co1233;
    full_adder adder1233(k12_33, co1233, k11_33, A[12] & B[21], co1232);
    wire k12_34;
    wire co1234;
    full_adder adder1234(k12_34, co1234, k11_34, A[12] & B[22], co1233);
    wire k12_35;
    wire co1235;
    full_adder adder1235(k12_35, co1235, k11_35, A[12] & B[23], co1234);
    wire k12_36;
    wire co1236;
    full_adder adder1236(k12_36, co1236, k11_36, A[12] & B[24], co1235);
    wire k12_37;
    wire co1237;
    full_adder adder1237(k12_37, co1237, k11_37, A[12] & B[25], co1236);
    wire k12_38;
    wire co1238;
    full_adder adder1238(k12_38, co1238, k11_38, A[12] & B[26], co1237);
    wire k12_39;
    wire co1239;
    full_adder adder1239(k12_39, co1239, k11_39, A[12] & B[27], co1238);
    wire k12_40;
    wire co1240;
    full_adder adder1240(k12_40, co1240, k11_40, A[12] & B[28], co1239);
    wire k12_41;
    wire co1241;
    full_adder adder1241(k12_41, co1241, k11_41, A[12] & B[29], co1240);
    wire k12_42;
    wire co1242;
    full_adder adder1242(k12_42, co1242, k11_42, A[12] & B[30], co1241);
    wire k12_43;
    wire co1243;
    full_adder adder1243(k12_43, co1243, co1142, !(A[12] & B[31]), co1242);
    // Row 13
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k13_13;
    wire co1313;
    full_adder adder1313(k13_13, co1313, k12_13, A[13] & B[0], 1'b0);
    wire k13_14;
    wire co1314;
    full_adder adder1314(k13_14, co1314, k12_14, A[13] & B[1], co1313);
    wire k13_15;
    wire co1315;
    full_adder adder1315(k13_15, co1315, k12_15, A[13] & B[2], co1314);
    wire k13_16;
    wire co1316;
    full_adder adder1316(k13_16, co1316, k12_16, A[13] & B[3], co1315);
    wire k13_17;
    wire co1317;
    full_adder adder1317(k13_17, co1317, k12_17, A[13] & B[4], co1316);
    wire k13_18;
    wire co1318;
    full_adder adder1318(k13_18, co1318, k12_18, A[13] & B[5], co1317);
    wire k13_19;
    wire co1319;
    full_adder adder1319(k13_19, co1319, k12_19, A[13] & B[6], co1318);
    wire k13_20;
    wire co1320;
    full_adder adder1320(k13_20, co1320, k12_20, A[13] & B[7], co1319);
    wire k13_21;
    wire co1321;
    full_adder adder1321(k13_21, co1321, k12_21, A[13] & B[8], co1320);
    wire k13_22;
    wire co1322;
    full_adder adder1322(k13_22, co1322, k12_22, A[13] & B[9], co1321);
    wire k13_23;
    wire co1323;
    full_adder adder1323(k13_23, co1323, k12_23, A[13] & B[10], co1322);
    wire k13_24;
    wire co1324;
    full_adder adder1324(k13_24, co1324, k12_24, A[13] & B[11], co1323);
    wire k13_25;
    wire co1325;
    full_adder adder1325(k13_25, co1325, k12_25, A[13] & B[12], co1324);
    wire k13_26;
    wire co1326;
    full_adder adder1326(k13_26, co1326, k12_26, A[13] & B[13], co1325);
    wire k13_27;
    wire co1327;
    full_adder adder1327(k13_27, co1327, k12_27, A[13] & B[14], co1326);
    wire k13_28;
    wire co1328;
    full_adder adder1328(k13_28, co1328, k12_28, A[13] & B[15], co1327);
    wire k13_29;
    wire co1329;
    full_adder adder1329(k13_29, co1329, k12_29, A[13] & B[16], co1328);
    wire k13_30;
    wire co1330;
    full_adder adder1330(k13_30, co1330, k12_30, A[13] & B[17], co1329);
    wire k13_31;
    wire co1331;
    full_adder adder1331(k13_31, co1331, k12_31, A[13] & B[18], co1330);
    wire k13_32;
    wire co1332;
    full_adder adder1332(k13_32, co1332, k12_32, A[13] & B[19], co1331);
    wire k13_33;
    wire co1333;
    full_adder adder1333(k13_33, co1333, k12_33, A[13] & B[20], co1332);
    wire k13_34;
    wire co1334;
    full_adder adder1334(k13_34, co1334, k12_34, A[13] & B[21], co1333);
    wire k13_35;
    wire co1335;
    full_adder adder1335(k13_35, co1335, k12_35, A[13] & B[22], co1334);
    wire k13_36;
    wire co1336;
    full_adder adder1336(k13_36, co1336, k12_36, A[13] & B[23], co1335);
    wire k13_37;
    wire co1337;
    full_adder adder1337(k13_37, co1337, k12_37, A[13] & B[24], co1336);
    wire k13_38;
    wire co1338;
    full_adder adder1338(k13_38, co1338, k12_38, A[13] & B[25], co1337);
    wire k13_39;
    wire co1339;
    full_adder adder1339(k13_39, co1339, k12_39, A[13] & B[26], co1338);
    wire k13_40;
    wire co1340;
    full_adder adder1340(k13_40, co1340, k12_40, A[13] & B[27], co1339);
    wire k13_41;
    wire co1341;
    full_adder adder1341(k13_41, co1341, k12_41, A[13] & B[28], co1340);
    wire k13_42;
    wire co1342;
    full_adder adder1342(k13_42, co1342, k12_42, A[13] & B[29], co1341);
    wire k13_43;
    wire co1343;
    full_adder adder1343(k13_43, co1343, k12_43, A[13] & B[30], co1342);
    wire k13_44;
    wire co1344;
    full_adder adder1344(k13_44, co1344, co1243, !(A[13] & B[31]), co1343);
    // Row 14
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k14_14;
    wire co1414;
    full_adder adder1414(k14_14, co1414, k13_14, A[14] & B[0], 1'b0);
    wire k14_15;
    wire co1415;
    full_adder adder1415(k14_15, co1415, k13_15, A[14] & B[1], co1414);
    wire k14_16;
    wire co1416;
    full_adder adder1416(k14_16, co1416, k13_16, A[14] & B[2], co1415);
    wire k14_17;
    wire co1417;
    full_adder adder1417(k14_17, co1417, k13_17, A[14] & B[3], co1416);
    wire k14_18;
    wire co1418;
    full_adder adder1418(k14_18, co1418, k13_18, A[14] & B[4], co1417);
    wire k14_19;
    wire co1419;
    full_adder adder1419(k14_19, co1419, k13_19, A[14] & B[5], co1418);
    wire k14_20;
    wire co1420;
    full_adder adder1420(k14_20, co1420, k13_20, A[14] & B[6], co1419);
    wire k14_21;
    wire co1421;
    full_adder adder1421(k14_21, co1421, k13_21, A[14] & B[7], co1420);
    wire k14_22;
    wire co1422;
    full_adder adder1422(k14_22, co1422, k13_22, A[14] & B[8], co1421);
    wire k14_23;
    wire co1423;
    full_adder adder1423(k14_23, co1423, k13_23, A[14] & B[9], co1422);
    wire k14_24;
    wire co1424;
    full_adder adder1424(k14_24, co1424, k13_24, A[14] & B[10], co1423);
    wire k14_25;
    wire co1425;
    full_adder adder1425(k14_25, co1425, k13_25, A[14] & B[11], co1424);
    wire k14_26;
    wire co1426;
    full_adder adder1426(k14_26, co1426, k13_26, A[14] & B[12], co1425);
    wire k14_27;
    wire co1427;
    full_adder adder1427(k14_27, co1427, k13_27, A[14] & B[13], co1426);
    wire k14_28;
    wire co1428;
    full_adder adder1428(k14_28, co1428, k13_28, A[14] & B[14], co1427);
    wire k14_29;
    wire co1429;
    full_adder adder1429(k14_29, co1429, k13_29, A[14] & B[15], co1428);
    wire k14_30;
    wire co1430;
    full_adder adder1430(k14_30, co1430, k13_30, A[14] & B[16], co1429);
    wire k14_31;
    wire co1431;
    full_adder adder1431(k14_31, co1431, k13_31, A[14] & B[17], co1430);
    wire k14_32;
    wire co1432;
    full_adder adder1432(k14_32, co1432, k13_32, A[14] & B[18], co1431);
    wire k14_33;
    wire co1433;
    full_adder adder1433(k14_33, co1433, k13_33, A[14] & B[19], co1432);
    wire k14_34;
    wire co1434;
    full_adder adder1434(k14_34, co1434, k13_34, A[14] & B[20], co1433);
    wire k14_35;
    wire co1435;
    full_adder adder1435(k14_35, co1435, k13_35, A[14] & B[21], co1434);
    wire k14_36;
    wire co1436;
    full_adder adder1436(k14_36, co1436, k13_36, A[14] & B[22], co1435);
    wire k14_37;
    wire co1437;
    full_adder adder1437(k14_37, co1437, k13_37, A[14] & B[23], co1436);
    wire k14_38;
    wire co1438;
    full_adder adder1438(k14_38, co1438, k13_38, A[14] & B[24], co1437);
    wire k14_39;
    wire co1439;
    full_adder adder1439(k14_39, co1439, k13_39, A[14] & B[25], co1438);
    wire k14_40;
    wire co1440;
    full_adder adder1440(k14_40, co1440, k13_40, A[14] & B[26], co1439);
    wire k14_41;
    wire co1441;
    full_adder adder1441(k14_41, co1441, k13_41, A[14] & B[27], co1440);
    wire k14_42;
    wire co1442;
    full_adder adder1442(k14_42, co1442, k13_42, A[14] & B[28], co1441);
    wire k14_43;
    wire co1443;
    full_adder adder1443(k14_43, co1443, k13_43, A[14] & B[29], co1442);
    wire k14_44;
    wire co1444;
    full_adder adder1444(k14_44, co1444, k13_44, A[14] & B[30], co1443);
    wire k14_45;
    wire co1445;
    full_adder adder1445(k14_45, co1445, co1344, !(A[14] & B[31]), co1444);
    // Row 15
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k15_15;
    wire co1515;
    full_adder adder1515(k15_15, co1515, k14_15, A[15] & B[0], 1'b0);
    wire k15_16;
    wire co1516;
    full_adder adder1516(k15_16, co1516, k14_16, A[15] & B[1], co1515);
    wire k15_17;
    wire co1517;
    full_adder adder1517(k15_17, co1517, k14_17, A[15] & B[2], co1516);
    wire k15_18;
    wire co1518;
    full_adder adder1518(k15_18, co1518, k14_18, A[15] & B[3], co1517);
    wire k15_19;
    wire co1519;
    full_adder adder1519(k15_19, co1519, k14_19, A[15] & B[4], co1518);
    wire k15_20;
    wire co1520;
    full_adder adder1520(k15_20, co1520, k14_20, A[15] & B[5], co1519);
    wire k15_21;
    wire co1521;
    full_adder adder1521(k15_21, co1521, k14_21, A[15] & B[6], co1520);
    wire k15_22;
    wire co1522;
    full_adder adder1522(k15_22, co1522, k14_22, A[15] & B[7], co1521);
    wire k15_23;
    wire co1523;
    full_adder adder1523(k15_23, co1523, k14_23, A[15] & B[8], co1522);
    wire k15_24;
    wire co1524;
    full_adder adder1524(k15_24, co1524, k14_24, A[15] & B[9], co1523);
    wire k15_25;
    wire co1525;
    full_adder adder1525(k15_25, co1525, k14_25, A[15] & B[10], co1524);
    wire k15_26;
    wire co1526;
    full_adder adder1526(k15_26, co1526, k14_26, A[15] & B[11], co1525);
    wire k15_27;
    wire co1527;
    full_adder adder1527(k15_27, co1527, k14_27, A[15] & B[12], co1526);
    wire k15_28;
    wire co1528;
    full_adder adder1528(k15_28, co1528, k14_28, A[15] & B[13], co1527);
    wire k15_29;
    wire co1529;
    full_adder adder1529(k15_29, co1529, k14_29, A[15] & B[14], co1528);
    wire k15_30;
    wire co1530;
    full_adder adder1530(k15_30, co1530, k14_30, A[15] & B[15], co1529);
    wire k15_31;
    wire co1531;
    full_adder adder1531(k15_31, co1531, k14_31, A[15] & B[16], co1530);
    wire k15_32;
    wire co1532;
    full_adder adder1532(k15_32, co1532, k14_32, A[15] & B[17], co1531);
    wire k15_33;
    wire co1533;
    full_adder adder1533(k15_33, co1533, k14_33, A[15] & B[18], co1532);
    wire k15_34;
    wire co1534;
    full_adder adder1534(k15_34, co1534, k14_34, A[15] & B[19], co1533);
    wire k15_35;
    wire co1535;
    full_adder adder1535(k15_35, co1535, k14_35, A[15] & B[20], co1534);
    wire k15_36;
    wire co1536;
    full_adder adder1536(k15_36, co1536, k14_36, A[15] & B[21], co1535);
    wire k15_37;
    wire co1537;
    full_adder adder1537(k15_37, co1537, k14_37, A[15] & B[22], co1536);
    wire k15_38;
    wire co1538;
    full_adder adder1538(k15_38, co1538, k14_38, A[15] & B[23], co1537);
    wire k15_39;
    wire co1539;
    full_adder adder1539(k15_39, co1539, k14_39, A[15] & B[24], co1538);
    wire k15_40;
    wire co1540;
    full_adder adder1540(k15_40, co1540, k14_40, A[15] & B[25], co1539);
    wire k15_41;
    wire co1541;
    full_adder adder1541(k15_41, co1541, k14_41, A[15] & B[26], co1540);
    wire k15_42;
    wire co1542;
    full_adder adder1542(k15_42, co1542, k14_42, A[15] & B[27], co1541);
    wire k15_43;
    wire co1543;
    full_adder adder1543(k15_43, co1543, k14_43, A[15] & B[28], co1542);
    wire k15_44;
    wire co1544;
    full_adder adder1544(k15_44, co1544, k14_44, A[15] & B[29], co1543);
    wire k15_45;
    wire co1545;
    full_adder adder1545(k15_45, co1545, k14_45, A[15] & B[30], co1544);
    wire k15_46;
    wire co1546;
    full_adder adder1546(k15_46, co1546, co1445, !(A[15] & B[31]), co1545);
    // Row 16
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k16_16;
    wire co1616;
    full_adder adder1616(k16_16, co1616, k15_16, A[16] & B[0], 1'b0);
    wire k16_17;
    wire co1617;
    full_adder adder1617(k16_17, co1617, k15_17, A[16] & B[1], co1616);
    wire k16_18;
    wire co1618;
    full_adder adder1618(k16_18, co1618, k15_18, A[16] & B[2], co1617);
    wire k16_19;
    wire co1619;
    full_adder adder1619(k16_19, co1619, k15_19, A[16] & B[3], co1618);
    wire k16_20;
    wire co1620;
    full_adder adder1620(k16_20, co1620, k15_20, A[16] & B[4], co1619);
    wire k16_21;
    wire co1621;
    full_adder adder1621(k16_21, co1621, k15_21, A[16] & B[5], co1620);
    wire k16_22;
    wire co1622;
    full_adder adder1622(k16_22, co1622, k15_22, A[16] & B[6], co1621);
    wire k16_23;
    wire co1623;
    full_adder adder1623(k16_23, co1623, k15_23, A[16] & B[7], co1622);
    wire k16_24;
    wire co1624;
    full_adder adder1624(k16_24, co1624, k15_24, A[16] & B[8], co1623);
    wire k16_25;
    wire co1625;
    full_adder adder1625(k16_25, co1625, k15_25, A[16] & B[9], co1624);
    wire k16_26;
    wire co1626;
    full_adder adder1626(k16_26, co1626, k15_26, A[16] & B[10], co1625);
    wire k16_27;
    wire co1627;
    full_adder adder1627(k16_27, co1627, k15_27, A[16] & B[11], co1626);
    wire k16_28;
    wire co1628;
    full_adder adder1628(k16_28, co1628, k15_28, A[16] & B[12], co1627);
    wire k16_29;
    wire co1629;
    full_adder adder1629(k16_29, co1629, k15_29, A[16] & B[13], co1628);
    wire k16_30;
    wire co1630;
    full_adder adder1630(k16_30, co1630, k15_30, A[16] & B[14], co1629);
    wire k16_31;
    wire co1631;
    full_adder adder1631(k16_31, co1631, k15_31, A[16] & B[15], co1630);
    wire k16_32;
    wire co1632;
    full_adder adder1632(k16_32, co1632, k15_32, A[16] & B[16], co1631);
    wire k16_33;
    wire co1633;
    full_adder adder1633(k16_33, co1633, k15_33, A[16] & B[17], co1632);
    wire k16_34;
    wire co1634;
    full_adder adder1634(k16_34, co1634, k15_34, A[16] & B[18], co1633);
    wire k16_35;
    wire co1635;
    full_adder adder1635(k16_35, co1635, k15_35, A[16] & B[19], co1634);
    wire k16_36;
    wire co1636;
    full_adder adder1636(k16_36, co1636, k15_36, A[16] & B[20], co1635);
    wire k16_37;
    wire co1637;
    full_adder adder1637(k16_37, co1637, k15_37, A[16] & B[21], co1636);
    wire k16_38;
    wire co1638;
    full_adder adder1638(k16_38, co1638, k15_38, A[16] & B[22], co1637);
    wire k16_39;
    wire co1639;
    full_adder adder1639(k16_39, co1639, k15_39, A[16] & B[23], co1638);
    wire k16_40;
    wire co1640;
    full_adder adder1640(k16_40, co1640, k15_40, A[16] & B[24], co1639);
    wire k16_41;
    wire co1641;
    full_adder adder1641(k16_41, co1641, k15_41, A[16] & B[25], co1640);
    wire k16_42;
    wire co1642;
    full_adder adder1642(k16_42, co1642, k15_42, A[16] & B[26], co1641);
    wire k16_43;
    wire co1643;
    full_adder adder1643(k16_43, co1643, k15_43, A[16] & B[27], co1642);
    wire k16_44;
    wire co1644;
    full_adder adder1644(k16_44, co1644, k15_44, A[16] & B[28], co1643);
    wire k16_45;
    wire co1645;
    full_adder adder1645(k16_45, co1645, k15_45, A[16] & B[29], co1644);
    wire k16_46;
    wire co1646;
    full_adder adder1646(k16_46, co1646, k15_46, A[16] & B[30], co1645);
    wire k16_47;
    wire co1647;
    full_adder adder1647(k16_47, co1647, co1546, !(A[16] & B[31]), co1646);
    // Row 17
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k17_17;
    wire co1717;
    full_adder adder1717(k17_17, co1717, k16_17, A[17] & B[0], 1'b0);
    wire k17_18;
    wire co1718;
    full_adder adder1718(k17_18, co1718, k16_18, A[17] & B[1], co1717);
    wire k17_19;
    wire co1719;
    full_adder adder1719(k17_19, co1719, k16_19, A[17] & B[2], co1718);
    wire k17_20;
    wire co1720;
    full_adder adder1720(k17_20, co1720, k16_20, A[17] & B[3], co1719);
    wire k17_21;
    wire co1721;
    full_adder adder1721(k17_21, co1721, k16_21, A[17] & B[4], co1720);
    wire k17_22;
    wire co1722;
    full_adder adder1722(k17_22, co1722, k16_22, A[17] & B[5], co1721);
    wire k17_23;
    wire co1723;
    full_adder adder1723(k17_23, co1723, k16_23, A[17] & B[6], co1722);
    wire k17_24;
    wire co1724;
    full_adder adder1724(k17_24, co1724, k16_24, A[17] & B[7], co1723);
    wire k17_25;
    wire co1725;
    full_adder adder1725(k17_25, co1725, k16_25, A[17] & B[8], co1724);
    wire k17_26;
    wire co1726;
    full_adder adder1726(k17_26, co1726, k16_26, A[17] & B[9], co1725);
    wire k17_27;
    wire co1727;
    full_adder adder1727(k17_27, co1727, k16_27, A[17] & B[10], co1726);
    wire k17_28;
    wire co1728;
    full_adder adder1728(k17_28, co1728, k16_28, A[17] & B[11], co1727);
    wire k17_29;
    wire co1729;
    full_adder adder1729(k17_29, co1729, k16_29, A[17] & B[12], co1728);
    wire k17_30;
    wire co1730;
    full_adder adder1730(k17_30, co1730, k16_30, A[17] & B[13], co1729);
    wire k17_31;
    wire co1731;
    full_adder adder1731(k17_31, co1731, k16_31, A[17] & B[14], co1730);
    wire k17_32;
    wire co1732;
    full_adder adder1732(k17_32, co1732, k16_32, A[17] & B[15], co1731);
    wire k17_33;
    wire co1733;
    full_adder adder1733(k17_33, co1733, k16_33, A[17] & B[16], co1732);
    wire k17_34;
    wire co1734;
    full_adder adder1734(k17_34, co1734, k16_34, A[17] & B[17], co1733);
    wire k17_35;
    wire co1735;
    full_adder adder1735(k17_35, co1735, k16_35, A[17] & B[18], co1734);
    wire k17_36;
    wire co1736;
    full_adder adder1736(k17_36, co1736, k16_36, A[17] & B[19], co1735);
    wire k17_37;
    wire co1737;
    full_adder adder1737(k17_37, co1737, k16_37, A[17] & B[20], co1736);
    wire k17_38;
    wire co1738;
    full_adder adder1738(k17_38, co1738, k16_38, A[17] & B[21], co1737);
    wire k17_39;
    wire co1739;
    full_adder adder1739(k17_39, co1739, k16_39, A[17] & B[22], co1738);
    wire k17_40;
    wire co1740;
    full_adder adder1740(k17_40, co1740, k16_40, A[17] & B[23], co1739);
    wire k17_41;
    wire co1741;
    full_adder adder1741(k17_41, co1741, k16_41, A[17] & B[24], co1740);
    wire k17_42;
    wire co1742;
    full_adder adder1742(k17_42, co1742, k16_42, A[17] & B[25], co1741);
    wire k17_43;
    wire co1743;
    full_adder adder1743(k17_43, co1743, k16_43, A[17] & B[26], co1742);
    wire k17_44;
    wire co1744;
    full_adder adder1744(k17_44, co1744, k16_44, A[17] & B[27], co1743);
    wire k17_45;
    wire co1745;
    full_adder adder1745(k17_45, co1745, k16_45, A[17] & B[28], co1744);
    wire k17_46;
    wire co1746;
    full_adder adder1746(k17_46, co1746, k16_46, A[17] & B[29], co1745);
    wire k17_47;
    wire co1747;
    full_adder adder1747(k17_47, co1747, k16_47, A[17] & B[30], co1746);
    wire k17_48;
    wire co1748;
    full_adder adder1748(k17_48, co1748, co1647, !(A[17] & B[31]), co1747);
    // Row 18
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k18_18;
    wire co1818;
    full_adder adder1818(k18_18, co1818, k17_18, A[18] & B[0], 1'b0);
    wire k18_19;
    wire co1819;
    full_adder adder1819(k18_19, co1819, k17_19, A[18] & B[1], co1818);
    wire k18_20;
    wire co1820;
    full_adder adder1820(k18_20, co1820, k17_20, A[18] & B[2], co1819);
    wire k18_21;
    wire co1821;
    full_adder adder1821(k18_21, co1821, k17_21, A[18] & B[3], co1820);
    wire k18_22;
    wire co1822;
    full_adder adder1822(k18_22, co1822, k17_22, A[18] & B[4], co1821);
    wire k18_23;
    wire co1823;
    full_adder adder1823(k18_23, co1823, k17_23, A[18] & B[5], co1822);
    wire k18_24;
    wire co1824;
    full_adder adder1824(k18_24, co1824, k17_24, A[18] & B[6], co1823);
    wire k18_25;
    wire co1825;
    full_adder adder1825(k18_25, co1825, k17_25, A[18] & B[7], co1824);
    wire k18_26;
    wire co1826;
    full_adder adder1826(k18_26, co1826, k17_26, A[18] & B[8], co1825);
    wire k18_27;
    wire co1827;
    full_adder adder1827(k18_27, co1827, k17_27, A[18] & B[9], co1826);
    wire k18_28;
    wire co1828;
    full_adder adder1828(k18_28, co1828, k17_28, A[18] & B[10], co1827);
    wire k18_29;
    wire co1829;
    full_adder adder1829(k18_29, co1829, k17_29, A[18] & B[11], co1828);
    wire k18_30;
    wire co1830;
    full_adder adder1830(k18_30, co1830, k17_30, A[18] & B[12], co1829);
    wire k18_31;
    wire co1831;
    full_adder adder1831(k18_31, co1831, k17_31, A[18] & B[13], co1830);
    wire k18_32;
    wire co1832;
    full_adder adder1832(k18_32, co1832, k17_32, A[18] & B[14], co1831);
    wire k18_33;
    wire co1833;
    full_adder adder1833(k18_33, co1833, k17_33, A[18] & B[15], co1832);
    wire k18_34;
    wire co1834;
    full_adder adder1834(k18_34, co1834, k17_34, A[18] & B[16], co1833);
    wire k18_35;
    wire co1835;
    full_adder adder1835(k18_35, co1835, k17_35, A[18] & B[17], co1834);
    wire k18_36;
    wire co1836;
    full_adder adder1836(k18_36, co1836, k17_36, A[18] & B[18], co1835);
    wire k18_37;
    wire co1837;
    full_adder adder1837(k18_37, co1837, k17_37, A[18] & B[19], co1836);
    wire k18_38;
    wire co1838;
    full_adder adder1838(k18_38, co1838, k17_38, A[18] & B[20], co1837);
    wire k18_39;
    wire co1839;
    full_adder adder1839(k18_39, co1839, k17_39, A[18] & B[21], co1838);
    wire k18_40;
    wire co1840;
    full_adder adder1840(k18_40, co1840, k17_40, A[18] & B[22], co1839);
    wire k18_41;
    wire co1841;
    full_adder adder1841(k18_41, co1841, k17_41, A[18] & B[23], co1840);
    wire k18_42;
    wire co1842;
    full_adder adder1842(k18_42, co1842, k17_42, A[18] & B[24], co1841);
    wire k18_43;
    wire co1843;
    full_adder adder1843(k18_43, co1843, k17_43, A[18] & B[25], co1842);
    wire k18_44;
    wire co1844;
    full_adder adder1844(k18_44, co1844, k17_44, A[18] & B[26], co1843);
    wire k18_45;
    wire co1845;
    full_adder adder1845(k18_45, co1845, k17_45, A[18] & B[27], co1844);
    wire k18_46;
    wire co1846;
    full_adder adder1846(k18_46, co1846, k17_46, A[18] & B[28], co1845);
    wire k18_47;
    wire co1847;
    full_adder adder1847(k18_47, co1847, k17_47, A[18] & B[29], co1846);
    wire k18_48;
    wire co1848;
    full_adder adder1848(k18_48, co1848, k17_48, A[18] & B[30], co1847);
    wire k18_49;
    wire co1849;
    full_adder adder1849(k18_49, co1849, co1748, !(A[18] & B[31]), co1848);
    // Row 19
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k19_19;
    wire co1919;
    full_adder adder1919(k19_19, co1919, k18_19, A[19] & B[0], 1'b0);
    wire k19_20;
    wire co1920;
    full_adder adder1920(k19_20, co1920, k18_20, A[19] & B[1], co1919);
    wire k19_21;
    wire co1921;
    full_adder adder1921(k19_21, co1921, k18_21, A[19] & B[2], co1920);
    wire k19_22;
    wire co1922;
    full_adder adder1922(k19_22, co1922, k18_22, A[19] & B[3], co1921);
    wire k19_23;
    wire co1923;
    full_adder adder1923(k19_23, co1923, k18_23, A[19] & B[4], co1922);
    wire k19_24;
    wire co1924;
    full_adder adder1924(k19_24, co1924, k18_24, A[19] & B[5], co1923);
    wire k19_25;
    wire co1925;
    full_adder adder1925(k19_25, co1925, k18_25, A[19] & B[6], co1924);
    wire k19_26;
    wire co1926;
    full_adder adder1926(k19_26, co1926, k18_26, A[19] & B[7], co1925);
    wire k19_27;
    wire co1927;
    full_adder adder1927(k19_27, co1927, k18_27, A[19] & B[8], co1926);
    wire k19_28;
    wire co1928;
    full_adder adder1928(k19_28, co1928, k18_28, A[19] & B[9], co1927);
    wire k19_29;
    wire co1929;
    full_adder adder1929(k19_29, co1929, k18_29, A[19] & B[10], co1928);
    wire k19_30;
    wire co1930;
    full_adder adder1930(k19_30, co1930, k18_30, A[19] & B[11], co1929);
    wire k19_31;
    wire co1931;
    full_adder adder1931(k19_31, co1931, k18_31, A[19] & B[12], co1930);
    wire k19_32;
    wire co1932;
    full_adder adder1932(k19_32, co1932, k18_32, A[19] & B[13], co1931);
    wire k19_33;
    wire co1933;
    full_adder adder1933(k19_33, co1933, k18_33, A[19] & B[14], co1932);
    wire k19_34;
    wire co1934;
    full_adder adder1934(k19_34, co1934, k18_34, A[19] & B[15], co1933);
    wire k19_35;
    wire co1935;
    full_adder adder1935(k19_35, co1935, k18_35, A[19] & B[16], co1934);
    wire k19_36;
    wire co1936;
    full_adder adder1936(k19_36, co1936, k18_36, A[19] & B[17], co1935);
    wire k19_37;
    wire co1937;
    full_adder adder1937(k19_37, co1937, k18_37, A[19] & B[18], co1936);
    wire k19_38;
    wire co1938;
    full_adder adder1938(k19_38, co1938, k18_38, A[19] & B[19], co1937);
    wire k19_39;
    wire co1939;
    full_adder adder1939(k19_39, co1939, k18_39, A[19] & B[20], co1938);
    wire k19_40;
    wire co1940;
    full_adder adder1940(k19_40, co1940, k18_40, A[19] & B[21], co1939);
    wire k19_41;
    wire co1941;
    full_adder adder1941(k19_41, co1941, k18_41, A[19] & B[22], co1940);
    wire k19_42;
    wire co1942;
    full_adder adder1942(k19_42, co1942, k18_42, A[19] & B[23], co1941);
    wire k19_43;
    wire co1943;
    full_adder adder1943(k19_43, co1943, k18_43, A[19] & B[24], co1942);
    wire k19_44;
    wire co1944;
    full_adder adder1944(k19_44, co1944, k18_44, A[19] & B[25], co1943);
    wire k19_45;
    wire co1945;
    full_adder adder1945(k19_45, co1945, k18_45, A[19] & B[26], co1944);
    wire k19_46;
    wire co1946;
    full_adder adder1946(k19_46, co1946, k18_46, A[19] & B[27], co1945);
    wire k19_47;
    wire co1947;
    full_adder adder1947(k19_47, co1947, k18_47, A[19] & B[28], co1946);
    wire k19_48;
    wire co1948;
    full_adder adder1948(k19_48, co1948, k18_48, A[19] & B[29], co1947);
    wire k19_49;
    wire co1949;
    full_adder adder1949(k19_49, co1949, k18_49, A[19] & B[30], co1948);
    wire k19_50;
    wire co1950;
    full_adder adder1950(k19_50, co1950, co1849, !(A[19] & B[31]), co1949);
    // Row 20
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k20_20;
    wire co2020;
    full_adder adder2020(k20_20, co2020, k19_20, A[20] & B[0], 1'b0);
    wire k20_21;
    wire co2021;
    full_adder adder2021(k20_21, co2021, k19_21, A[20] & B[1], co2020);
    wire k20_22;
    wire co2022;
    full_adder adder2022(k20_22, co2022, k19_22, A[20] & B[2], co2021);
    wire k20_23;
    wire co2023;
    full_adder adder2023(k20_23, co2023, k19_23, A[20] & B[3], co2022);
    wire k20_24;
    wire co2024;
    full_adder adder2024(k20_24, co2024, k19_24, A[20] & B[4], co2023);
    wire k20_25;
    wire co2025;
    full_adder adder2025(k20_25, co2025, k19_25, A[20] & B[5], co2024);
    wire k20_26;
    wire co2026;
    full_adder adder2026(k20_26, co2026, k19_26, A[20] & B[6], co2025);
    wire k20_27;
    wire co2027;
    full_adder adder2027(k20_27, co2027, k19_27, A[20] & B[7], co2026);
    wire k20_28;
    wire co2028;
    full_adder adder2028(k20_28, co2028, k19_28, A[20] & B[8], co2027);
    wire k20_29;
    wire co2029;
    full_adder adder2029(k20_29, co2029, k19_29, A[20] & B[9], co2028);
    wire k20_30;
    wire co2030;
    full_adder adder2030(k20_30, co2030, k19_30, A[20] & B[10], co2029);
    wire k20_31;
    wire co2031;
    full_adder adder2031(k20_31, co2031, k19_31, A[20] & B[11], co2030);
    wire k20_32;
    wire co2032;
    full_adder adder2032(k20_32, co2032, k19_32, A[20] & B[12], co2031);
    wire k20_33;
    wire co2033;
    full_adder adder2033(k20_33, co2033, k19_33, A[20] & B[13], co2032);
    wire k20_34;
    wire co2034;
    full_adder adder2034(k20_34, co2034, k19_34, A[20] & B[14], co2033);
    wire k20_35;
    wire co2035;
    full_adder adder2035(k20_35, co2035, k19_35, A[20] & B[15], co2034);
    wire k20_36;
    wire co2036;
    full_adder adder2036(k20_36, co2036, k19_36, A[20] & B[16], co2035);
    wire k20_37;
    wire co2037;
    full_adder adder2037(k20_37, co2037, k19_37, A[20] & B[17], co2036);
    wire k20_38;
    wire co2038;
    full_adder adder2038(k20_38, co2038, k19_38, A[20] & B[18], co2037);
    wire k20_39;
    wire co2039;
    full_adder adder2039(k20_39, co2039, k19_39, A[20] & B[19], co2038);
    wire k20_40;
    wire co2040;
    full_adder adder2040(k20_40, co2040, k19_40, A[20] & B[20], co2039);
    wire k20_41;
    wire co2041;
    full_adder adder2041(k20_41, co2041, k19_41, A[20] & B[21], co2040);
    wire k20_42;
    wire co2042;
    full_adder adder2042(k20_42, co2042, k19_42, A[20] & B[22], co2041);
    wire k20_43;
    wire co2043;
    full_adder adder2043(k20_43, co2043, k19_43, A[20] & B[23], co2042);
    wire k20_44;
    wire co2044;
    full_adder adder2044(k20_44, co2044, k19_44, A[20] & B[24], co2043);
    wire k20_45;
    wire co2045;
    full_adder adder2045(k20_45, co2045, k19_45, A[20] & B[25], co2044);
    wire k20_46;
    wire co2046;
    full_adder adder2046(k20_46, co2046, k19_46, A[20] & B[26], co2045);
    wire k20_47;
    wire co2047;
    full_adder adder2047(k20_47, co2047, k19_47, A[20] & B[27], co2046);
    wire k20_48;
    wire co2048;
    full_adder adder2048(k20_48, co2048, k19_48, A[20] & B[28], co2047);
    wire k20_49;
    wire co2049;
    full_adder adder2049(k20_49, co2049, k19_49, A[20] & B[29], co2048);
    wire k20_50;
    wire co2050;
    full_adder adder2050(k20_50, co2050, k19_50, A[20] & B[30], co2049);
    wire k20_51;
    wire co2051;
    full_adder adder2051(k20_51, co2051, co1950, !(A[20] & B[31]), co2050);
    // Row 21
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k21_21;
    wire co2121;
    full_adder adder2121(k21_21, co2121, k20_21, A[21] & B[0], 1'b0);
    wire k21_22;
    wire co2122;
    full_adder adder2122(k21_22, co2122, k20_22, A[21] & B[1], co2121);
    wire k21_23;
    wire co2123;
    full_adder adder2123(k21_23, co2123, k20_23, A[21] & B[2], co2122);
    wire k21_24;
    wire co2124;
    full_adder adder2124(k21_24, co2124, k20_24, A[21] & B[3], co2123);
    wire k21_25;
    wire co2125;
    full_adder adder2125(k21_25, co2125, k20_25, A[21] & B[4], co2124);
    wire k21_26;
    wire co2126;
    full_adder adder2126(k21_26, co2126, k20_26, A[21] & B[5], co2125);
    wire k21_27;
    wire co2127;
    full_adder adder2127(k21_27, co2127, k20_27, A[21] & B[6], co2126);
    wire k21_28;
    wire co2128;
    full_adder adder2128(k21_28, co2128, k20_28, A[21] & B[7], co2127);
    wire k21_29;
    wire co2129;
    full_adder adder2129(k21_29, co2129, k20_29, A[21] & B[8], co2128);
    wire k21_30;
    wire co2130;
    full_adder adder2130(k21_30, co2130, k20_30, A[21] & B[9], co2129);
    wire k21_31;
    wire co2131;
    full_adder adder2131(k21_31, co2131, k20_31, A[21] & B[10], co2130);
    wire k21_32;
    wire co2132;
    full_adder adder2132(k21_32, co2132, k20_32, A[21] & B[11], co2131);
    wire k21_33;
    wire co2133;
    full_adder adder2133(k21_33, co2133, k20_33, A[21] & B[12], co2132);
    wire k21_34;
    wire co2134;
    full_adder adder2134(k21_34, co2134, k20_34, A[21] & B[13], co2133);
    wire k21_35;
    wire co2135;
    full_adder adder2135(k21_35, co2135, k20_35, A[21] & B[14], co2134);
    wire k21_36;
    wire co2136;
    full_adder adder2136(k21_36, co2136, k20_36, A[21] & B[15], co2135);
    wire k21_37;
    wire co2137;
    full_adder adder2137(k21_37, co2137, k20_37, A[21] & B[16], co2136);
    wire k21_38;
    wire co2138;
    full_adder adder2138(k21_38, co2138, k20_38, A[21] & B[17], co2137);
    wire k21_39;
    wire co2139;
    full_adder adder2139(k21_39, co2139, k20_39, A[21] & B[18], co2138);
    wire k21_40;
    wire co2140;
    full_adder adder2140(k21_40, co2140, k20_40, A[21] & B[19], co2139);
    wire k21_41;
    wire co2141;
    full_adder adder2141(k21_41, co2141, k20_41, A[21] & B[20], co2140);
    wire k21_42;
    wire co2142;
    full_adder adder2142(k21_42, co2142, k20_42, A[21] & B[21], co2141);
    wire k21_43;
    wire co2143;
    full_adder adder2143(k21_43, co2143, k20_43, A[21] & B[22], co2142);
    wire k21_44;
    wire co2144;
    full_adder adder2144(k21_44, co2144, k20_44, A[21] & B[23], co2143);
    wire k21_45;
    wire co2145;
    full_adder adder2145(k21_45, co2145, k20_45, A[21] & B[24], co2144);
    wire k21_46;
    wire co2146;
    full_adder adder2146(k21_46, co2146, k20_46, A[21] & B[25], co2145);
    wire k21_47;
    wire co2147;
    full_adder adder2147(k21_47, co2147, k20_47, A[21] & B[26], co2146);
    wire k21_48;
    wire co2148;
    full_adder adder2148(k21_48, co2148, k20_48, A[21] & B[27], co2147);
    wire k21_49;
    wire co2149;
    full_adder adder2149(k21_49, co2149, k20_49, A[21] & B[28], co2148);
    wire k21_50;
    wire co2150;
    full_adder adder2150(k21_50, co2150, k20_50, A[21] & B[29], co2149);
    wire k21_51;
    wire co2151;
    full_adder adder2151(k21_51, co2151, k20_51, A[21] & B[30], co2150);
    wire k21_52;
    wire co2152;
    full_adder adder2152(k21_52, co2152, co2051, !(A[21] & B[31]), co2151);
    // Row 22
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k22_22;
    wire co2222;
    full_adder adder2222(k22_22, co2222, k21_22, A[22] & B[0], 1'b0);
    wire k22_23;
    wire co2223;
    full_adder adder2223(k22_23, co2223, k21_23, A[22] & B[1], co2222);
    wire k22_24;
    wire co2224;
    full_adder adder2224(k22_24, co2224, k21_24, A[22] & B[2], co2223);
    wire k22_25;
    wire co2225;
    full_adder adder2225(k22_25, co2225, k21_25, A[22] & B[3], co2224);
    wire k22_26;
    wire co2226;
    full_adder adder2226(k22_26, co2226, k21_26, A[22] & B[4], co2225);
    wire k22_27;
    wire co2227;
    full_adder adder2227(k22_27, co2227, k21_27, A[22] & B[5], co2226);
    wire k22_28;
    wire co2228;
    full_adder adder2228(k22_28, co2228, k21_28, A[22] & B[6], co2227);
    wire k22_29;
    wire co2229;
    full_adder adder2229(k22_29, co2229, k21_29, A[22] & B[7], co2228);
    wire k22_30;
    wire co2230;
    full_adder adder2230(k22_30, co2230, k21_30, A[22] & B[8], co2229);
    wire k22_31;
    wire co2231;
    full_adder adder2231(k22_31, co2231, k21_31, A[22] & B[9], co2230);
    wire k22_32;
    wire co2232;
    full_adder adder2232(k22_32, co2232, k21_32, A[22] & B[10], co2231);
    wire k22_33;
    wire co2233;
    full_adder adder2233(k22_33, co2233, k21_33, A[22] & B[11], co2232);
    wire k22_34;
    wire co2234;
    full_adder adder2234(k22_34, co2234, k21_34, A[22] & B[12], co2233);
    wire k22_35;
    wire co2235;
    full_adder adder2235(k22_35, co2235, k21_35, A[22] & B[13], co2234);
    wire k22_36;
    wire co2236;
    full_adder adder2236(k22_36, co2236, k21_36, A[22] & B[14], co2235);
    wire k22_37;
    wire co2237;
    full_adder adder2237(k22_37, co2237, k21_37, A[22] & B[15], co2236);
    wire k22_38;
    wire co2238;
    full_adder adder2238(k22_38, co2238, k21_38, A[22] & B[16], co2237);
    wire k22_39;
    wire co2239;
    full_adder adder2239(k22_39, co2239, k21_39, A[22] & B[17], co2238);
    wire k22_40;
    wire co2240;
    full_adder adder2240(k22_40, co2240, k21_40, A[22] & B[18], co2239);
    wire k22_41;
    wire co2241;
    full_adder adder2241(k22_41, co2241, k21_41, A[22] & B[19], co2240);
    wire k22_42;
    wire co2242;
    full_adder adder2242(k22_42, co2242, k21_42, A[22] & B[20], co2241);
    wire k22_43;
    wire co2243;
    full_adder adder2243(k22_43, co2243, k21_43, A[22] & B[21], co2242);
    wire k22_44;
    wire co2244;
    full_adder adder2244(k22_44, co2244, k21_44, A[22] & B[22], co2243);
    wire k22_45;
    wire co2245;
    full_adder adder2245(k22_45, co2245, k21_45, A[22] & B[23], co2244);
    wire k22_46;
    wire co2246;
    full_adder adder2246(k22_46, co2246, k21_46, A[22] & B[24], co2245);
    wire k22_47;
    wire co2247;
    full_adder adder2247(k22_47, co2247, k21_47, A[22] & B[25], co2246);
    wire k22_48;
    wire co2248;
    full_adder adder2248(k22_48, co2248, k21_48, A[22] & B[26], co2247);
    wire k22_49;
    wire co2249;
    full_adder adder2249(k22_49, co2249, k21_49, A[22] & B[27], co2248);
    wire k22_50;
    wire co2250;
    full_adder adder2250(k22_50, co2250, k21_50, A[22] & B[28], co2249);
    wire k22_51;
    wire co2251;
    full_adder adder2251(k22_51, co2251, k21_51, A[22] & B[29], co2250);
    wire k22_52;
    wire co2252;
    full_adder adder2252(k22_52, co2252, k21_52, A[22] & B[30], co2251);
    wire k22_53;
    wire co2253;
    full_adder adder2253(k22_53, co2253, co2152, !(A[22] & B[31]), co2252);
    // Row 23
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k23_23;
    wire co2323;
    full_adder adder2323(k23_23, co2323, k22_23, A[23] & B[0], 1'b0);
    wire k23_24;
    wire co2324;
    full_adder adder2324(k23_24, co2324, k22_24, A[23] & B[1], co2323);
    wire k23_25;
    wire co2325;
    full_adder adder2325(k23_25, co2325, k22_25, A[23] & B[2], co2324);
    wire k23_26;
    wire co2326;
    full_adder adder2326(k23_26, co2326, k22_26, A[23] & B[3], co2325);
    wire k23_27;
    wire co2327;
    full_adder adder2327(k23_27, co2327, k22_27, A[23] & B[4], co2326);
    wire k23_28;
    wire co2328;
    full_adder adder2328(k23_28, co2328, k22_28, A[23] & B[5], co2327);
    wire k23_29;
    wire co2329;
    full_adder adder2329(k23_29, co2329, k22_29, A[23] & B[6], co2328);
    wire k23_30;
    wire co2330;
    full_adder adder2330(k23_30, co2330, k22_30, A[23] & B[7], co2329);
    wire k23_31;
    wire co2331;
    full_adder adder2331(k23_31, co2331, k22_31, A[23] & B[8], co2330);
    wire k23_32;
    wire co2332;
    full_adder adder2332(k23_32, co2332, k22_32, A[23] & B[9], co2331);
    wire k23_33;
    wire co2333;
    full_adder adder2333(k23_33, co2333, k22_33, A[23] & B[10], co2332);
    wire k23_34;
    wire co2334;
    full_adder adder2334(k23_34, co2334, k22_34, A[23] & B[11], co2333);
    wire k23_35;
    wire co2335;
    full_adder adder2335(k23_35, co2335, k22_35, A[23] & B[12], co2334);
    wire k23_36;
    wire co2336;
    full_adder adder2336(k23_36, co2336, k22_36, A[23] & B[13], co2335);
    wire k23_37;
    wire co2337;
    full_adder adder2337(k23_37, co2337, k22_37, A[23] & B[14], co2336);
    wire k23_38;
    wire co2338;
    full_adder adder2338(k23_38, co2338, k22_38, A[23] & B[15], co2337);
    wire k23_39;
    wire co2339;
    full_adder adder2339(k23_39, co2339, k22_39, A[23] & B[16], co2338);
    wire k23_40;
    wire co2340;
    full_adder adder2340(k23_40, co2340, k22_40, A[23] & B[17], co2339);
    wire k23_41;
    wire co2341;
    full_adder adder2341(k23_41, co2341, k22_41, A[23] & B[18], co2340);
    wire k23_42;
    wire co2342;
    full_adder adder2342(k23_42, co2342, k22_42, A[23] & B[19], co2341);
    wire k23_43;
    wire co2343;
    full_adder adder2343(k23_43, co2343, k22_43, A[23] & B[20], co2342);
    wire k23_44;
    wire co2344;
    full_adder adder2344(k23_44, co2344, k22_44, A[23] & B[21], co2343);
    wire k23_45;
    wire co2345;
    full_adder adder2345(k23_45, co2345, k22_45, A[23] & B[22], co2344);
    wire k23_46;
    wire co2346;
    full_adder adder2346(k23_46, co2346, k22_46, A[23] & B[23], co2345);
    wire k23_47;
    wire co2347;
    full_adder adder2347(k23_47, co2347, k22_47, A[23] & B[24], co2346);
    wire k23_48;
    wire co2348;
    full_adder adder2348(k23_48, co2348, k22_48, A[23] & B[25], co2347);
    wire k23_49;
    wire co2349;
    full_adder adder2349(k23_49, co2349, k22_49, A[23] & B[26], co2348);
    wire k23_50;
    wire co2350;
    full_adder adder2350(k23_50, co2350, k22_50, A[23] & B[27], co2349);
    wire k23_51;
    wire co2351;
    full_adder adder2351(k23_51, co2351, k22_51, A[23] & B[28], co2350);
    wire k23_52;
    wire co2352;
    full_adder adder2352(k23_52, co2352, k22_52, A[23] & B[29], co2351);
    wire k23_53;
    wire co2353;
    full_adder adder2353(k23_53, co2353, k22_53, A[23] & B[30], co2352);
    wire k23_54;
    wire co2354;
    full_adder adder2354(k23_54, co2354, co2253, !(A[23] & B[31]), co2353);
    // Row 24
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k24_24;
    wire co2424;
    full_adder adder2424(k24_24, co2424, k23_24, A[24] & B[0], 1'b0);
    wire k24_25;
    wire co2425;
    full_adder adder2425(k24_25, co2425, k23_25, A[24] & B[1], co2424);
    wire k24_26;
    wire co2426;
    full_adder adder2426(k24_26, co2426, k23_26, A[24] & B[2], co2425);
    wire k24_27;
    wire co2427;
    full_adder adder2427(k24_27, co2427, k23_27, A[24] & B[3], co2426);
    wire k24_28;
    wire co2428;
    full_adder adder2428(k24_28, co2428, k23_28, A[24] & B[4], co2427);
    wire k24_29;
    wire co2429;
    full_adder adder2429(k24_29, co2429, k23_29, A[24] & B[5], co2428);
    wire k24_30;
    wire co2430;
    full_adder adder2430(k24_30, co2430, k23_30, A[24] & B[6], co2429);
    wire k24_31;
    wire co2431;
    full_adder adder2431(k24_31, co2431, k23_31, A[24] & B[7], co2430);
    wire k24_32;
    wire co2432;
    full_adder adder2432(k24_32, co2432, k23_32, A[24] & B[8], co2431);
    wire k24_33;
    wire co2433;
    full_adder adder2433(k24_33, co2433, k23_33, A[24] & B[9], co2432);
    wire k24_34;
    wire co2434;
    full_adder adder2434(k24_34, co2434, k23_34, A[24] & B[10], co2433);
    wire k24_35;
    wire co2435;
    full_adder adder2435(k24_35, co2435, k23_35, A[24] & B[11], co2434);
    wire k24_36;
    wire co2436;
    full_adder adder2436(k24_36, co2436, k23_36, A[24] & B[12], co2435);
    wire k24_37;
    wire co2437;
    full_adder adder2437(k24_37, co2437, k23_37, A[24] & B[13], co2436);
    wire k24_38;
    wire co2438;
    full_adder adder2438(k24_38, co2438, k23_38, A[24] & B[14], co2437);
    wire k24_39;
    wire co2439;
    full_adder adder2439(k24_39, co2439, k23_39, A[24] & B[15], co2438);
    wire k24_40;
    wire co2440;
    full_adder adder2440(k24_40, co2440, k23_40, A[24] & B[16], co2439);
    wire k24_41;
    wire co2441;
    full_adder adder2441(k24_41, co2441, k23_41, A[24] & B[17], co2440);
    wire k24_42;
    wire co2442;
    full_adder adder2442(k24_42, co2442, k23_42, A[24] & B[18], co2441);
    wire k24_43;
    wire co2443;
    full_adder adder2443(k24_43, co2443, k23_43, A[24] & B[19], co2442);
    wire k24_44;
    wire co2444;
    full_adder adder2444(k24_44, co2444, k23_44, A[24] & B[20], co2443);
    wire k24_45;
    wire co2445;
    full_adder adder2445(k24_45, co2445, k23_45, A[24] & B[21], co2444);
    wire k24_46;
    wire co2446;
    full_adder adder2446(k24_46, co2446, k23_46, A[24] & B[22], co2445);
    wire k24_47;
    wire co2447;
    full_adder adder2447(k24_47, co2447, k23_47, A[24] & B[23], co2446);
    wire k24_48;
    wire co2448;
    full_adder adder2448(k24_48, co2448, k23_48, A[24] & B[24], co2447);
    wire k24_49;
    wire co2449;
    full_adder adder2449(k24_49, co2449, k23_49, A[24] & B[25], co2448);
    wire k24_50;
    wire co2450;
    full_adder adder2450(k24_50, co2450, k23_50, A[24] & B[26], co2449);
    wire k24_51;
    wire co2451;
    full_adder adder2451(k24_51, co2451, k23_51, A[24] & B[27], co2450);
    wire k24_52;
    wire co2452;
    full_adder adder2452(k24_52, co2452, k23_52, A[24] & B[28], co2451);
    wire k24_53;
    wire co2453;
    full_adder adder2453(k24_53, co2453, k23_53, A[24] & B[29], co2452);
    wire k24_54;
    wire co2454;
    full_adder adder2454(k24_54, co2454, k23_54, A[24] & B[30], co2453);
    wire k24_55;
    wire co2455;
    full_adder adder2455(k24_55, co2455, co2354, !(A[24] & B[31]), co2454);
    // Row 25
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k25_25;
    wire co2525;
    full_adder adder2525(k25_25, co2525, k24_25, A[25] & B[0], 1'b0);
    wire k25_26;
    wire co2526;
    full_adder adder2526(k25_26, co2526, k24_26, A[25] & B[1], co2525);
    wire k25_27;
    wire co2527;
    full_adder adder2527(k25_27, co2527, k24_27, A[25] & B[2], co2526);
    wire k25_28;
    wire co2528;
    full_adder adder2528(k25_28, co2528, k24_28, A[25] & B[3], co2527);
    wire k25_29;
    wire co2529;
    full_adder adder2529(k25_29, co2529, k24_29, A[25] & B[4], co2528);
    wire k25_30;
    wire co2530;
    full_adder adder2530(k25_30, co2530, k24_30, A[25] & B[5], co2529);
    wire k25_31;
    wire co2531;
    full_adder adder2531(k25_31, co2531, k24_31, A[25] & B[6], co2530);
    wire k25_32;
    wire co2532;
    full_adder adder2532(k25_32, co2532, k24_32, A[25] & B[7], co2531);
    wire k25_33;
    wire co2533;
    full_adder adder2533(k25_33, co2533, k24_33, A[25] & B[8], co2532);
    wire k25_34;
    wire co2534;
    full_adder adder2534(k25_34, co2534, k24_34, A[25] & B[9], co2533);
    wire k25_35;
    wire co2535;
    full_adder adder2535(k25_35, co2535, k24_35, A[25] & B[10], co2534);
    wire k25_36;
    wire co2536;
    full_adder adder2536(k25_36, co2536, k24_36, A[25] & B[11], co2535);
    wire k25_37;
    wire co2537;
    full_adder adder2537(k25_37, co2537, k24_37, A[25] & B[12], co2536);
    wire k25_38;
    wire co2538;
    full_adder adder2538(k25_38, co2538, k24_38, A[25] & B[13], co2537);
    wire k25_39;
    wire co2539;
    full_adder adder2539(k25_39, co2539, k24_39, A[25] & B[14], co2538);
    wire k25_40;
    wire co2540;
    full_adder adder2540(k25_40, co2540, k24_40, A[25] & B[15], co2539);
    wire k25_41;
    wire co2541;
    full_adder adder2541(k25_41, co2541, k24_41, A[25] & B[16], co2540);
    wire k25_42;
    wire co2542;
    full_adder adder2542(k25_42, co2542, k24_42, A[25] & B[17], co2541);
    wire k25_43;
    wire co2543;
    full_adder adder2543(k25_43, co2543, k24_43, A[25] & B[18], co2542);
    wire k25_44;
    wire co2544;
    full_adder adder2544(k25_44, co2544, k24_44, A[25] & B[19], co2543);
    wire k25_45;
    wire co2545;
    full_adder adder2545(k25_45, co2545, k24_45, A[25] & B[20], co2544);
    wire k25_46;
    wire co2546;
    full_adder adder2546(k25_46, co2546, k24_46, A[25] & B[21], co2545);
    wire k25_47;
    wire co2547;
    full_adder adder2547(k25_47, co2547, k24_47, A[25] & B[22], co2546);
    wire k25_48;
    wire co2548;
    full_adder adder2548(k25_48, co2548, k24_48, A[25] & B[23], co2547);
    wire k25_49;
    wire co2549;
    full_adder adder2549(k25_49, co2549, k24_49, A[25] & B[24], co2548);
    wire k25_50;
    wire co2550;
    full_adder adder2550(k25_50, co2550, k24_50, A[25] & B[25], co2549);
    wire k25_51;
    wire co2551;
    full_adder adder2551(k25_51, co2551, k24_51, A[25] & B[26], co2550);
    wire k25_52;
    wire co2552;
    full_adder adder2552(k25_52, co2552, k24_52, A[25] & B[27], co2551);
    wire k25_53;
    wire co2553;
    full_adder adder2553(k25_53, co2553, k24_53, A[25] & B[28], co2552);
    wire k25_54;
    wire co2554;
    full_adder adder2554(k25_54, co2554, k24_54, A[25] & B[29], co2553);
    wire k25_55;
    wire co2555;
    full_adder adder2555(k25_55, co2555, k24_55, A[25] & B[30], co2554);
    wire k25_56;
    wire co2556;
    full_adder adder2556(k25_56, co2556, co2455, !(A[25] & B[31]), co2555);
    // Row 26
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k26_26;
    wire co2626;
    full_adder adder2626(k26_26, co2626, k25_26, A[26] & B[0], 1'b0);
    wire k26_27;
    wire co2627;
    full_adder adder2627(k26_27, co2627, k25_27, A[26] & B[1], co2626);
    wire k26_28;
    wire co2628;
    full_adder adder2628(k26_28, co2628, k25_28, A[26] & B[2], co2627);
    wire k26_29;
    wire co2629;
    full_adder adder2629(k26_29, co2629, k25_29, A[26] & B[3], co2628);
    wire k26_30;
    wire co2630;
    full_adder adder2630(k26_30, co2630, k25_30, A[26] & B[4], co2629);
    wire k26_31;
    wire co2631;
    full_adder adder2631(k26_31, co2631, k25_31, A[26] & B[5], co2630);
    wire k26_32;
    wire co2632;
    full_adder adder2632(k26_32, co2632, k25_32, A[26] & B[6], co2631);
    wire k26_33;
    wire co2633;
    full_adder adder2633(k26_33, co2633, k25_33, A[26] & B[7], co2632);
    wire k26_34;
    wire co2634;
    full_adder adder2634(k26_34, co2634, k25_34, A[26] & B[8], co2633);
    wire k26_35;
    wire co2635;
    full_adder adder2635(k26_35, co2635, k25_35, A[26] & B[9], co2634);
    wire k26_36;
    wire co2636;
    full_adder adder2636(k26_36, co2636, k25_36, A[26] & B[10], co2635);
    wire k26_37;
    wire co2637;
    full_adder adder2637(k26_37, co2637, k25_37, A[26] & B[11], co2636);
    wire k26_38;
    wire co2638;
    full_adder adder2638(k26_38, co2638, k25_38, A[26] & B[12], co2637);
    wire k26_39;
    wire co2639;
    full_adder adder2639(k26_39, co2639, k25_39, A[26] & B[13], co2638);
    wire k26_40;
    wire co2640;
    full_adder adder2640(k26_40, co2640, k25_40, A[26] & B[14], co2639);
    wire k26_41;
    wire co2641;
    full_adder adder2641(k26_41, co2641, k25_41, A[26] & B[15], co2640);
    wire k26_42;
    wire co2642;
    full_adder adder2642(k26_42, co2642, k25_42, A[26] & B[16], co2641);
    wire k26_43;
    wire co2643;
    full_adder adder2643(k26_43, co2643, k25_43, A[26] & B[17], co2642);
    wire k26_44;
    wire co2644;
    full_adder adder2644(k26_44, co2644, k25_44, A[26] & B[18], co2643);
    wire k26_45;
    wire co2645;
    full_adder adder2645(k26_45, co2645, k25_45, A[26] & B[19], co2644);
    wire k26_46;
    wire co2646;
    full_adder adder2646(k26_46, co2646, k25_46, A[26] & B[20], co2645);
    wire k26_47;
    wire co2647;
    full_adder adder2647(k26_47, co2647, k25_47, A[26] & B[21], co2646);
    wire k26_48;
    wire co2648;
    full_adder adder2648(k26_48, co2648, k25_48, A[26] & B[22], co2647);
    wire k26_49;
    wire co2649;
    full_adder adder2649(k26_49, co2649, k25_49, A[26] & B[23], co2648);
    wire k26_50;
    wire co2650;
    full_adder adder2650(k26_50, co2650, k25_50, A[26] & B[24], co2649);
    wire k26_51;
    wire co2651;
    full_adder adder2651(k26_51, co2651, k25_51, A[26] & B[25], co2650);
    wire k26_52;
    wire co2652;
    full_adder adder2652(k26_52, co2652, k25_52, A[26] & B[26], co2651);
    wire k26_53;
    wire co2653;
    full_adder adder2653(k26_53, co2653, k25_53, A[26] & B[27], co2652);
    wire k26_54;
    wire co2654;
    full_adder adder2654(k26_54, co2654, k25_54, A[26] & B[28], co2653);
    wire k26_55;
    wire co2655;
    full_adder adder2655(k26_55, co2655, k25_55, A[26] & B[29], co2654);
    wire k26_56;
    wire co2656;
    full_adder adder2656(k26_56, co2656, k25_56, A[26] & B[30], co2655);
    wire k26_57;
    wire co2657;
    full_adder adder2657(k26_57, co2657, co2556, !(A[26] & B[31]), co2656);
    // Row 27
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k27_27;
    wire co2727;
    full_adder adder2727(k27_27, co2727, k26_27, A[27] & B[0], 1'b0);
    wire k27_28;
    wire co2728;
    full_adder adder2728(k27_28, co2728, k26_28, A[27] & B[1], co2727);
    wire k27_29;
    wire co2729;
    full_adder adder2729(k27_29, co2729, k26_29, A[27] & B[2], co2728);
    wire k27_30;
    wire co2730;
    full_adder adder2730(k27_30, co2730, k26_30, A[27] & B[3], co2729);
    wire k27_31;
    wire co2731;
    full_adder adder2731(k27_31, co2731, k26_31, A[27] & B[4], co2730);
    wire k27_32;
    wire co2732;
    full_adder adder2732(k27_32, co2732, k26_32, A[27] & B[5], co2731);
    wire k27_33;
    wire co2733;
    full_adder adder2733(k27_33, co2733, k26_33, A[27] & B[6], co2732);
    wire k27_34;
    wire co2734;
    full_adder adder2734(k27_34, co2734, k26_34, A[27] & B[7], co2733);
    wire k27_35;
    wire co2735;
    full_adder adder2735(k27_35, co2735, k26_35, A[27] & B[8], co2734);
    wire k27_36;
    wire co2736;
    full_adder adder2736(k27_36, co2736, k26_36, A[27] & B[9], co2735);
    wire k27_37;
    wire co2737;
    full_adder adder2737(k27_37, co2737, k26_37, A[27] & B[10], co2736);
    wire k27_38;
    wire co2738;
    full_adder adder2738(k27_38, co2738, k26_38, A[27] & B[11], co2737);
    wire k27_39;
    wire co2739;
    full_adder adder2739(k27_39, co2739, k26_39, A[27] & B[12], co2738);
    wire k27_40;
    wire co2740;
    full_adder adder2740(k27_40, co2740, k26_40, A[27] & B[13], co2739);
    wire k27_41;
    wire co2741;
    full_adder adder2741(k27_41, co2741, k26_41, A[27] & B[14], co2740);
    wire k27_42;
    wire co2742;
    full_adder adder2742(k27_42, co2742, k26_42, A[27] & B[15], co2741);
    wire k27_43;
    wire co2743;
    full_adder adder2743(k27_43, co2743, k26_43, A[27] & B[16], co2742);
    wire k27_44;
    wire co2744;
    full_adder adder2744(k27_44, co2744, k26_44, A[27] & B[17], co2743);
    wire k27_45;
    wire co2745;
    full_adder adder2745(k27_45, co2745, k26_45, A[27] & B[18], co2744);
    wire k27_46;
    wire co2746;
    full_adder adder2746(k27_46, co2746, k26_46, A[27] & B[19], co2745);
    wire k27_47;
    wire co2747;
    full_adder adder2747(k27_47, co2747, k26_47, A[27] & B[20], co2746);
    wire k27_48;
    wire co2748;
    full_adder adder2748(k27_48, co2748, k26_48, A[27] & B[21], co2747);
    wire k27_49;
    wire co2749;
    full_adder adder2749(k27_49, co2749, k26_49, A[27] & B[22], co2748);
    wire k27_50;
    wire co2750;
    full_adder adder2750(k27_50, co2750, k26_50, A[27] & B[23], co2749);
    wire k27_51;
    wire co2751;
    full_adder adder2751(k27_51, co2751, k26_51, A[27] & B[24], co2750);
    wire k27_52;
    wire co2752;
    full_adder adder2752(k27_52, co2752, k26_52, A[27] & B[25], co2751);
    wire k27_53;
    wire co2753;
    full_adder adder2753(k27_53, co2753, k26_53, A[27] & B[26], co2752);
    wire k27_54;
    wire co2754;
    full_adder adder2754(k27_54, co2754, k26_54, A[27] & B[27], co2753);
    wire k27_55;
    wire co2755;
    full_adder adder2755(k27_55, co2755, k26_55, A[27] & B[28], co2754);
    wire k27_56;
    wire co2756;
    full_adder adder2756(k27_56, co2756, k26_56, A[27] & B[29], co2755);
    wire k27_57;
    wire co2757;
    full_adder adder2757(k27_57, co2757, k26_57, A[27] & B[30], co2756);
    wire k27_58;
    wire co2758;
    full_adder adder2758(k27_58, co2758, co2657, !(A[27] & B[31]), co2757);
    // Row 28
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k28_28;
    wire co2828;
    full_adder adder2828(k28_28, co2828, k27_28, A[28] & B[0], 1'b0);
    wire k28_29;
    wire co2829;
    full_adder adder2829(k28_29, co2829, k27_29, A[28] & B[1], co2828);
    wire k28_30;
    wire co2830;
    full_adder adder2830(k28_30, co2830, k27_30, A[28] & B[2], co2829);
    wire k28_31;
    wire co2831;
    full_adder adder2831(k28_31, co2831, k27_31, A[28] & B[3], co2830);
    wire k28_32;
    wire co2832;
    full_adder adder2832(k28_32, co2832, k27_32, A[28] & B[4], co2831);
    wire k28_33;
    wire co2833;
    full_adder adder2833(k28_33, co2833, k27_33, A[28] & B[5], co2832);
    wire k28_34;
    wire co2834;
    full_adder adder2834(k28_34, co2834, k27_34, A[28] & B[6], co2833);
    wire k28_35;
    wire co2835;
    full_adder adder2835(k28_35, co2835, k27_35, A[28] & B[7], co2834);
    wire k28_36;
    wire co2836;
    full_adder adder2836(k28_36, co2836, k27_36, A[28] & B[8], co2835);
    wire k28_37;
    wire co2837;
    full_adder adder2837(k28_37, co2837, k27_37, A[28] & B[9], co2836);
    wire k28_38;
    wire co2838;
    full_adder adder2838(k28_38, co2838, k27_38, A[28] & B[10], co2837);
    wire k28_39;
    wire co2839;
    full_adder adder2839(k28_39, co2839, k27_39, A[28] & B[11], co2838);
    wire k28_40;
    wire co2840;
    full_adder adder2840(k28_40, co2840, k27_40, A[28] & B[12], co2839);
    wire k28_41;
    wire co2841;
    full_adder adder2841(k28_41, co2841, k27_41, A[28] & B[13], co2840);
    wire k28_42;
    wire co2842;
    full_adder adder2842(k28_42, co2842, k27_42, A[28] & B[14], co2841);
    wire k28_43;
    wire co2843;
    full_adder adder2843(k28_43, co2843, k27_43, A[28] & B[15], co2842);
    wire k28_44;
    wire co2844;
    full_adder adder2844(k28_44, co2844, k27_44, A[28] & B[16], co2843);
    wire k28_45;
    wire co2845;
    full_adder adder2845(k28_45, co2845, k27_45, A[28] & B[17], co2844);
    wire k28_46;
    wire co2846;
    full_adder adder2846(k28_46, co2846, k27_46, A[28] & B[18], co2845);
    wire k28_47;
    wire co2847;
    full_adder adder2847(k28_47, co2847, k27_47, A[28] & B[19], co2846);
    wire k28_48;
    wire co2848;
    full_adder adder2848(k28_48, co2848, k27_48, A[28] & B[20], co2847);
    wire k28_49;
    wire co2849;
    full_adder adder2849(k28_49, co2849, k27_49, A[28] & B[21], co2848);
    wire k28_50;
    wire co2850;
    full_adder adder2850(k28_50, co2850, k27_50, A[28] & B[22], co2849);
    wire k28_51;
    wire co2851;
    full_adder adder2851(k28_51, co2851, k27_51, A[28] & B[23], co2850);
    wire k28_52;
    wire co2852;
    full_adder adder2852(k28_52, co2852, k27_52, A[28] & B[24], co2851);
    wire k28_53;
    wire co2853;
    full_adder adder2853(k28_53, co2853, k27_53, A[28] & B[25], co2852);
    wire k28_54;
    wire co2854;
    full_adder adder2854(k28_54, co2854, k27_54, A[28] & B[26], co2853);
    wire k28_55;
    wire co2855;
    full_adder adder2855(k28_55, co2855, k27_55, A[28] & B[27], co2854);
    wire k28_56;
    wire co2856;
    full_adder adder2856(k28_56, co2856, k27_56, A[28] & B[28], co2855);
    wire k28_57;
    wire co2857;
    full_adder adder2857(k28_57, co2857, k27_57, A[28] & B[29], co2856);
    wire k28_58;
    wire co2858;
    full_adder adder2858(k28_58, co2858, k27_58, A[28] & B[30], co2857);
    wire k28_59;
    wire co2859;
    full_adder adder2859(k28_59, co2859, co2758, !(A[28] & B[31]), co2858);
    // Row 29
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k29_29;
    wire co2929;
    full_adder adder2929(k29_29, co2929, k28_29, A[29] & B[0], 1'b0);
    wire k29_30;
    wire co2930;
    full_adder adder2930(k29_30, co2930, k28_30, A[29] & B[1], co2929);
    wire k29_31;
    wire co2931;
    full_adder adder2931(k29_31, co2931, k28_31, A[29] & B[2], co2930);
    wire k29_32;
    wire co2932;
    full_adder adder2932(k29_32, co2932, k28_32, A[29] & B[3], co2931);
    wire k29_33;
    wire co2933;
    full_adder adder2933(k29_33, co2933, k28_33, A[29] & B[4], co2932);
    wire k29_34;
    wire co2934;
    full_adder adder2934(k29_34, co2934, k28_34, A[29] & B[5], co2933);
    wire k29_35;
    wire co2935;
    full_adder adder2935(k29_35, co2935, k28_35, A[29] & B[6], co2934);
    wire k29_36;
    wire co2936;
    full_adder adder2936(k29_36, co2936, k28_36, A[29] & B[7], co2935);
    wire k29_37;
    wire co2937;
    full_adder adder2937(k29_37, co2937, k28_37, A[29] & B[8], co2936);
    wire k29_38;
    wire co2938;
    full_adder adder2938(k29_38, co2938, k28_38, A[29] & B[9], co2937);
    wire k29_39;
    wire co2939;
    full_adder adder2939(k29_39, co2939, k28_39, A[29] & B[10], co2938);
    wire k29_40;
    wire co2940;
    full_adder adder2940(k29_40, co2940, k28_40, A[29] & B[11], co2939);
    wire k29_41;
    wire co2941;
    full_adder adder2941(k29_41, co2941, k28_41, A[29] & B[12], co2940);
    wire k29_42;
    wire co2942;
    full_adder adder2942(k29_42, co2942, k28_42, A[29] & B[13], co2941);
    wire k29_43;
    wire co2943;
    full_adder adder2943(k29_43, co2943, k28_43, A[29] & B[14], co2942);
    wire k29_44;
    wire co2944;
    full_adder adder2944(k29_44, co2944, k28_44, A[29] & B[15], co2943);
    wire k29_45;
    wire co2945;
    full_adder adder2945(k29_45, co2945, k28_45, A[29] & B[16], co2944);
    wire k29_46;
    wire co2946;
    full_adder adder2946(k29_46, co2946, k28_46, A[29] & B[17], co2945);
    wire k29_47;
    wire co2947;
    full_adder adder2947(k29_47, co2947, k28_47, A[29] & B[18], co2946);
    wire k29_48;
    wire co2948;
    full_adder adder2948(k29_48, co2948, k28_48, A[29] & B[19], co2947);
    wire k29_49;
    wire co2949;
    full_adder adder2949(k29_49, co2949, k28_49, A[29] & B[20], co2948);
    wire k29_50;
    wire co2950;
    full_adder adder2950(k29_50, co2950, k28_50, A[29] & B[21], co2949);
    wire k29_51;
    wire co2951;
    full_adder adder2951(k29_51, co2951, k28_51, A[29] & B[22], co2950);
    wire k29_52;
    wire co2952;
    full_adder adder2952(k29_52, co2952, k28_52, A[29] & B[23], co2951);
    wire k29_53;
    wire co2953;
    full_adder adder2953(k29_53, co2953, k28_53, A[29] & B[24], co2952);
    wire k29_54;
    wire co2954;
    full_adder adder2954(k29_54, co2954, k28_54, A[29] & B[25], co2953);
    wire k29_55;
    wire co2955;
    full_adder adder2955(k29_55, co2955, k28_55, A[29] & B[26], co2954);
    wire k29_56;
    wire co2956;
    full_adder adder2956(k29_56, co2956, k28_56, A[29] & B[27], co2955);
    wire k29_57;
    wire co2957;
    full_adder adder2957(k29_57, co2957, k28_57, A[29] & B[28], co2956);
    wire k29_58;
    wire co2958;
    full_adder adder2958(k29_58, co2958, k28_58, A[29] & B[29], co2957);
    wire k29_59;
    wire co2959;
    full_adder adder2959(k29_59, co2959, k28_59, A[29] & B[30], co2958);
    wire k29_60;
    wire co2960;
    full_adder adder2960(k29_60, co2960, co2859, !(A[29] & B[31]), co2959);
    // Row 30
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k30_30;
    wire co3030;
    full_adder adder3030(k30_30, co3030, k29_30, A[30] & B[0], 1'b0);
    wire k30_31;
    wire co3031;
    full_adder adder3031(k30_31, co3031, k29_31, A[30] & B[1], co3030);
    wire k30_32;
    wire co3032;
    full_adder adder3032(k30_32, co3032, k29_32, A[30] & B[2], co3031);
    wire k30_33;
    wire co3033;
    full_adder adder3033(k30_33, co3033, k29_33, A[30] & B[3], co3032);
    wire k30_34;
    wire co3034;
    full_adder adder3034(k30_34, co3034, k29_34, A[30] & B[4], co3033);
    wire k30_35;
    wire co3035;
    full_adder adder3035(k30_35, co3035, k29_35, A[30] & B[5], co3034);
    wire k30_36;
    wire co3036;
    full_adder adder3036(k30_36, co3036, k29_36, A[30] & B[6], co3035);
    wire k30_37;
    wire co3037;
    full_adder adder3037(k30_37, co3037, k29_37, A[30] & B[7], co3036);
    wire k30_38;
    wire co3038;
    full_adder adder3038(k30_38, co3038, k29_38, A[30] & B[8], co3037);
    wire k30_39;
    wire co3039;
    full_adder adder3039(k30_39, co3039, k29_39, A[30] & B[9], co3038);
    wire k30_40;
    wire co3040;
    full_adder adder3040(k30_40, co3040, k29_40, A[30] & B[10], co3039);
    wire k30_41;
    wire co3041;
    full_adder adder3041(k30_41, co3041, k29_41, A[30] & B[11], co3040);
    wire k30_42;
    wire co3042;
    full_adder adder3042(k30_42, co3042, k29_42, A[30] & B[12], co3041);
    wire k30_43;
    wire co3043;
    full_adder adder3043(k30_43, co3043, k29_43, A[30] & B[13], co3042);
    wire k30_44;
    wire co3044;
    full_adder adder3044(k30_44, co3044, k29_44, A[30] & B[14], co3043);
    wire k30_45;
    wire co3045;
    full_adder adder3045(k30_45, co3045, k29_45, A[30] & B[15], co3044);
    wire k30_46;
    wire co3046;
    full_adder adder3046(k30_46, co3046, k29_46, A[30] & B[16], co3045);
    wire k30_47;
    wire co3047;
    full_adder adder3047(k30_47, co3047, k29_47, A[30] & B[17], co3046);
    wire k30_48;
    wire co3048;
    full_adder adder3048(k30_48, co3048, k29_48, A[30] & B[18], co3047);
    wire k30_49;
    wire co3049;
    full_adder adder3049(k30_49, co3049, k29_49, A[30] & B[19], co3048);
    wire k30_50;
    wire co3050;
    full_adder adder3050(k30_50, co3050, k29_50, A[30] & B[20], co3049);
    wire k30_51;
    wire co3051;
    full_adder adder3051(k30_51, co3051, k29_51, A[30] & B[21], co3050);
    wire k30_52;
    wire co3052;
    full_adder adder3052(k30_52, co3052, k29_52, A[30] & B[22], co3051);
    wire k30_53;
    wire co3053;
    full_adder adder3053(k30_53, co3053, k29_53, A[30] & B[23], co3052);
    wire k30_54;
    wire co3054;
    full_adder adder3054(k30_54, co3054, k29_54, A[30] & B[24], co3053);
    wire k30_55;
    wire co3055;
    full_adder adder3055(k30_55, co3055, k29_55, A[30] & B[25], co3054);
    wire k30_56;
    wire co3056;
    full_adder adder3056(k30_56, co3056, k29_56, A[30] & B[26], co3055);
    wire k30_57;
    wire co3057;
    full_adder adder3057(k30_57, co3057, k29_57, A[30] & B[27], co3056);
    wire k30_58;
    wire co3058;
    full_adder adder3058(k30_58, co3058, k29_58, A[30] & B[28], co3057);
    wire k30_59;
    wire co3059;
    full_adder adder3059(k30_59, co3059, k29_59, A[30] & B[29], co3058);
    wire k30_60;
    wire co3060;
    full_adder adder3060(k30_60, co3060, k29_60, A[30] & B[30], co3059);
    wire k30_61;
    wire co3061;
    full_adder adder3061(k30_61, co3061, co2960, !(A[30] & B[31]), co3060);
    // Row 31
    // Wires with k are outputs of the adders
    // Wires with co are carry outs
    wire k31_31;
    wire co3131;
    full_adder adder3131(k31_31, co3131, k30_31, !(A[31] & B[0]), 1'b0);
    wire k31_32;
    wire co3132;
    full_adder adder3132(k31_32, co3132, k30_32, !(A[31] & B[1]), co3131);
    wire k31_33;
    wire co3133;
    full_adder adder3133(k31_33, co3133, k30_33, !(A[31] & B[2]), co3132);
    wire k31_34;
    wire co3134;
    full_adder adder3134(k31_34, co3134, k30_34, !(A[31] & B[3]), co3133);
    wire k31_35;
    wire co3135;
    full_adder adder3135(k31_35, co3135, k30_35, !(A[31] & B[4]), co3134);
    wire k31_36;
    wire co3136;
    full_adder adder3136(k31_36, co3136, k30_36, !(A[31] & B[5]), co3135);
    wire k31_37;
    wire co3137;
    full_adder adder3137(k31_37, co3137, k30_37, !(A[31] & B[6]), co3136);
    wire k31_38;
    wire co3138;
    full_adder adder3138(k31_38, co3138, k30_38, !(A[31] & B[7]), co3137);
    wire k31_39;
    wire co3139;
    full_adder adder3139(k31_39, co3139, k30_39, !(A[31] & B[8]), co3138);
    wire k31_40;
    wire co3140;
    full_adder adder3140(k31_40, co3140, k30_40, !(A[31] & B[9]), co3139);
    wire k31_41;
    wire co3141;
    full_adder adder3141(k31_41, co3141, k30_41, !(A[31] & B[10]), co3140);
    wire k31_42;
    wire co3142;
    full_adder adder3142(k31_42, co3142, k30_42, !(A[31] & B[11]), co3141);
    wire k31_43;
    wire co3143;
    full_adder adder3143(k31_43, co3143, k30_43, !(A[31] & B[12]), co3142);
    wire k31_44;
    wire co3144;
    full_adder adder3144(k31_44, co3144, k30_44, !(A[31] & B[13]), co3143);
    wire k31_45;
    wire co3145;
    full_adder adder3145(k31_45, co3145, k30_45, !(A[31] & B[14]), co3144);
    wire k31_46;
    wire co3146;
    full_adder adder3146(k31_46, co3146, k30_46, !(A[31] & B[15]), co3145);
    wire k31_47;
    wire co3147;
    full_adder adder3147(k31_47, co3147, k30_47, !(A[31] & B[16]), co3146);
    wire k31_48;
    wire co3148;
    full_adder adder3148(k31_48, co3148, k30_48, !(A[31] & B[17]), co3147);
    wire k31_49;
    wire co3149;
    full_adder adder3149(k31_49, co3149, k30_49, !(A[31] & B[18]), co3148);
    wire k31_50;
    wire co3150;
    full_adder adder3150(k31_50, co3150, k30_50, !(A[31] & B[19]), co3149);
    wire k31_51;
    wire co3151;
    full_adder adder3151(k31_51, co3151, k30_51, !(A[31] & B[20]), co3150);
    wire k31_52;
    wire co3152;
    full_adder adder3152(k31_52, co3152, k30_52, !(A[31] & B[21]), co3151);
    wire k31_53;
    wire co3153;
    full_adder adder3153(k31_53, co3153, k30_53, !(A[31] & B[22]), co3152);
    wire k31_54;
    wire co3154;
    full_adder adder3154(k31_54, co3154, k30_54, !(A[31] & B[23]), co3153);
    wire k31_55;
    wire co3155;
    full_adder adder3155(k31_55, co3155, k30_55, !(A[31] & B[24]), co3154);
    wire k31_56;
    wire co3156;
    full_adder adder3156(k31_56, co3156, k30_56, !(A[31] & B[25]), co3155);
    wire k31_57;
    wire co3157;
    full_adder adder3157(k31_57, co3157, k30_57, !(A[31] & B[26]), co3156);
    wire k31_58;
    wire co3158;
    full_adder adder3158(k31_58, co3158, k30_58, !(A[31] & B[27]), co3157);
    wire k31_59;
    wire co3159;
    full_adder adder3159(k31_59, co3159, k30_59, !(A[31] & B[28]), co3158);
    wire k31_60;
    wire co3160;
    full_adder adder3160(k31_60, co3160, k30_60, !(A[31] & B[29]), co3159);
    wire k31_61;
    wire co3161;
    full_adder adder3161(k31_61, co3161, k30_61, !(A[31] & B[30]), co3160);
    wire k31_62;
    wire co3162;
    full_adder adder3162(k31_62, co3162, co3061, (A[31] & B[31]), co3161);

    assign O[0]  = k0_0;
    assign O[1]  = k1_1;
    assign O[2]  = k2_2;
    assign O[3]  = k3_3;
    assign O[4]  = k4_4;
    assign O[5]  = k5_5;
    assign O[6]  = k6_6;
    assign O[7]  = k7_7;
    assign O[8]  = k8_8;
    assign O[9]  = k9_9;
    assign O[10] = k10_10;
    assign O[11] = k11_11;
    assign O[12] = k12_12;
    assign O[13] = k13_13;
    assign O[14] = k14_14;
    assign O[15] = k15_15;
    assign O[16] = k16_16;
    assign O[17] = k17_17;
    assign O[18] = k18_18;
    assign O[19] = k19_19;
    assign O[20] = k20_20;
    assign O[21] = k21_21;
    assign O[22] = k22_22;
    assign O[23] = k23_23;
    assign O[24] = k24_24;
    assign O[25] = k25_25;
    assign O[26] = k26_26;
    assign O[27] = k27_27;
    assign O[28] = k28_28;
    assign O[29] = k29_29;
    assign O[30] = k30_30;
    assign O[31] = k31_31;

    assign O[32] = k31_32;
    assign O[33] = k31_33;
    assign O[34] = k31_34;
    assign O[35] = k31_35;
    assign O[36] = k31_36;
    assign O[37] = k31_37;
    assign O[38] = k31_38;
    assign O[39] = k31_39;
    assign O[40] = k31_40;
    assign O[41] = k31_41;
    assign O[42] = k31_42;
    assign O[43] = k31_43;
    assign O[44] = k31_44;
    assign O[45] = k31_45;
    assign O[46] = k31_46;
    assign O[47] = k31_47;
    assign O[48] = k31_48;
    assign O[49] = k31_49;
    assign O[50] = k31_50;
    assign O[51] = k31_51;
    assign O[52] = k31_52;
    assign O[53] = k31_53;
    assign O[54] = k31_54;
    assign O[55] = k31_55;
    assign O[56] = k31_56;
    assign O[57] = k31_57;
    assign O[58] = k31_58;
    assign O[59] = k31_59;
    assign O[60] = k31_60;
    assign O[61] = k31_61;
    assign O[62] = k31_62;
    
    //full_adder(S, Cout, A, B, Cin);

    wire trash;

    full_adder LAST(O[63], trash, 1'b1, 1'b0, co3162);
    //assign O[63] = co3162;


    // if you OR bits [63:31] and you get 1, and if you AND all the bits and you get 0, then there is overflow
    // if you OR bits [63:31] and you get 0, and if you AND all the bits and you get 1, then there is overflow
    output overflow;
    wire anded, ored;
    assign anded = &O[63:31];
    assign ored = |O[63:31];

    xor ovf(overflow, anded, ored);

    output ready;
    input clk, ctrl_MULT;

    wire [5:0] count;

    counter counttttttt(clk, ctrl_MULT, count);
    assign ready = ~count[5] & ~count[4] & count[3] & ~count[2] & ~count[1] & ~count[0];


endmodule